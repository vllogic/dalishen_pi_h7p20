// ============================================================
// File Name: tx_dpram_768x32_emif.v
// IP core  : ethernet_mac_v2 
// Function : TX memory management
// ============================================================

module cme_ip_tx_dpram_768x32_emif_v3(
        clkw,
        cew,
        aw,
        dw,
        wr_ram_sel,

        clkr,
        cer,
        ar,
        qr,
        mti_rdy_i,
        rd_ram_sel
        );
//protect_encode_begin
`pragma protect begin_protected
`pragma protect version=1
`pragma protect data_block
joqvu!!!dmls<joqvu!!!dfs<joqvu!!!xs`sbn`tfm<joqvu!!!se`sbn`tfm<joqvu!!!nuj`sez`j<joqvu!!!\9;1^!bs<pvuqvu!!\42;1^!rs<!!!!joqvu!!!dmlx<joqvu!!!dfx<joqvu!!!\21;1^!bx<joqvu!!!\8;1^!!ex<xjsf!nuj`sez`j<xjsf!fnc`df`s1`w1<xjsf!fnc`df`s1`w2<xjsf!fnc`df`s2`w1<xjsf!fnc`df`s2`w2<xjsf!fnc`df`s3`w2<xjsf!fnc`df`s3`w1<sfh!!\8;1^!!ex`mpx<sfh!!!!!!!!!bs`9`t<xjsf!\26;1^!ex`jo<xjsf!\8;1^!!bx`ijhi<xjsf!\42;1^!rs`1<xjsf!\42;1^!rs`2<xjsf!\42;1^!rs`3<bttjho!rs!>!se`sbn`tfm!@!)bs`9`t!@!rs`3!;!rs`2*!;!)bs`9`t!@!rs`3!;!rs`1*<!bmxbzt!A)qptfehf!dmls*!cfhjojg)nuj`sez`j*!!!bs`9`t!=>!bs\9^<foebmxbzt!A)qptfehf!dmlx*!cfhjojg)dfx!'!)bx\1^**!!!ex`mpx!=>!ex<foebttjho!ex`jo!>!bx\1^!@!|ex-ex`mpx~!;!|ex-ex~<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s1`w2)
!/dmlx)dmlx*-
!/bx)bx\:;3^*-
!/dfx)fnc`df`s1`w2*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`1\42;27^*!!!!*<bttjho!fnc`df`s1`w2!>!)xs`sbn`tfm*!'!)bx\21^*!'!bx\2^!'!dfx<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s1`w1)
!/dmlx)dmlx*-
!/bx)bx\:;3^*-
!/dfx)fnc`df`s1`w1*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`1\26;1^*!!!!*<bttjho!fnc`df`s1`w1!>!)xs`sbn`tfm*!'!)bx\21^*!'!)bx\2^*!'!dfx<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s2`w2)
!/dmlx)dmlx*-
!/bx)bx\:;3^*-
!/dfx)fnc`df`s2`w2*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`2\42;27^*!!!!*<bttjho!fnc`df`s2`w2!>!xs`sbn`tfm!'!)bx\21^*!'!bx\2^!'!dfx<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s2`w1)
!/dmlx)dmlx*-
!/bx)bx\:;3^*-
!/dfx)fnc`df`s2`w1*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`2\26;1^*!!!!*<bttjho!fnc`df`s2`w1!>!xs`sbn`tfm!'!)bx\21^*!'!)bx\2^*!'!dfx<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s3`w2)
!/dmlx)dmlx*-
!/bx)bx`ijhi*-
!/dfx)fnc`df`s3`w2*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`3\42;27^*!!!!*<bttjho!bx`ijhi!>!xs`sbn`tfm!@!|2(c2-bx\9;3^~!;!|2(c1-bx\9;3^~<bttjho!fnc`df`s3`w2!>!bx\21^!'!bx\2^!'!dfx<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s3`w1)
!/dmlx)dmlx*-
!/bx)bx`ijhi*-
!/dfx)fnc`df`s3`w1*-
!/ex)ex`jo*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs*-
!/rs)rs`3\26;1^*!!!!*<bttjho!fnc`df`s3`w1!>!bx\21^!'!)bx\2^*!'!dfx<
`pragma protect end_protected
//protect_encode_end
endmodule


