//================================================================================
// Copyright (c) 2013 Capital-micro, Inc.(Beijing)  All rights reserved.
//
// Capital-micro, Inc.(Beijing) Confidential.
//
// No part of this code may be reproduced, distributed, transmitted,
// transcribed, stored in a retrieval system, or translated into any
// human or computer language, in any form or by any means, electronic,
// mechanical, magnetic, manual, or otherwise, without the express
// written permission of Capital-micro, Inc.
//
//================================================================================
// Module Description: Transmit and Receive Memory Control
// This module is used to implement:
// 1. Transmit DPRAM Control
// 2. Receive DPRAM Control
// 3. Interface with ethernet MAC core 
//================================================================================
// Revision History :
//     V1.0   2013-03-18  FPGA IP Grp, first created
//     V2.0   2014-04-25  FPGA IP Grp, support EMIF/AHB bus, modify TX/RX
//     memory management
//     V3.0   2014-12-18  FPGA IP Grp, add eth_mac_core_f_1k.v to support
//     1000M mode 
//================================================================================

module hme_ip_tr_mem_ctrl_ahb_v3 (
   clk_app_i,
   clk_tx_i,
   clk_rx_i,

   rst_clk_app_n,
   rst_clk_tx_n,
   rst_clk_rx_n,

   // MAC Transmit interface
   mti_val_o,          
   mti_data_o,
   mti_sof_o,
   mti_eof_o,
   mti_be_o,
   mti_discrc_o,
   mti_dispad_o,
   mti_flowctrl_o,
   mti_rdy_i,
   mti_txstatus_i,
   mti_txstatus_val_i,
   // MAC Receive interface
   mri_val_i,      
   mri_data_i,
   mri_be_i,
   mri_sof_i,
   mri_eof_i,
   mri_rxstatus_i,
   //interface with emif2mci   
   tx_mem_wr,
   tx_mem_wr_addr,
   tx_mem_wr_data,   
   tx_stat_val_o,
   tx_stat,
   tx_mem_0_clr,
   tx_mem_1_clr,
   
   tx_mem_rd_en,

   mci_ctrl,

   rx_mem_rd,
   rx_mem_frame_len,
   rx_mem_frame_status,
   rx_mem_rd_data,
   rcv_new_frame_en_rx,
   rcv_new_frame_en_clr_app,
   frame_rd_over_en_pedge
);
`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
JZKHfPuSqfAmjPVbVxhSKtUcvcjPj6+4QCp6QiFxv4nsP111dMWg4lZnLvWHxZMziq4ZnoWMa3GvTlkfyAx459JwXYUp9++mcX9h4iv0ELA73xF35/nLcT+Xn0raOA2RiqLC1DolMQLhhJGzN4NnSkXeaeOgmwY/bEh2w9tyWiE=
`pragma protect data_block
6so86mxGW2+3cYvx+h5Cenn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3meWNhyezaw/77O5iSYNXTW15EDKLY2O7EBys0fWCGOv
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgeresZfHLsBYUVq8xpnpR22oashAaUCSqF8I4058We6jYP400x1UJ84KzJr+mVGIrQGE
Nklp2V1qKrauRKLYzeP1GCMPOcex85fJ8k/1Wo2NUfZHmAoyYomKoWlQi7pnZJepPn7+5K1rKNzS5ax7RgSfBnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3tHsqwAY+pfLcLvDJr55dFkRHq30AKqda5FHm2PDhNKb6so86mxGW2+3cYvx+h5Cenn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3tEeI90e8DHEL3ECxtkWaPhZmzceFvZIW0xIbCvfxbRr2l3gn2b1cMxTddGyYFaSfx3EusWfl9U8IgE2SqAXK9mAi440WLBSRtiqNNGWN7gw
0doLoChOBeXdY4l4gm9qzvdc9IexOoh0u/kbObv9SjrmLG6xoEdk3W8tci1nShx7Hywaw13UT4aZhfbQ+ub2mWt7EjsNZWqHiyUTMtph61yayWn/1EJx2Em2c938CLfd
NRaSL/AfN+0zowmgyyM4Tf9NLANrtWzSx4z6iXJgziTcMxhyWTyhSP9wm7ID1uNUDnE3tr/6SNkCk+FRLVsjlpGsWswcVMZklAi5nQ7hJRWp4qs2wJUzcCxc4d7RST3s
C2ECLe5tHsZv3brOzlgylWAmpaqmeKqE20zzZUP8xtzuBTzI2j34NYnBJoAjm5I4CH4q/feIL6jQou/Ppwl65x95tl2wChGLWs/Akzr5MZVdzyZXG5+cgZxZIXcUTTg2
yh2LZBS/bPrQnH6yeS4vi5rJaf/UQnHYSbZz3fwIt936N3nvCIitArLzpx09/LXryWa8b0xgUnemYhdi/6PJpkzVCrbTvRrixTx4q0IwAQHcNi4K3jscbo1Jj4vhxqdd
mslp/9RCcdhJtnPd/Ai33bBAIFPBueWV5l37MZzWkzjjHspMoeXY7O1KrIKIF2IdvkaQpSShwLHfWhpVTpvBps+kI1RwRzLCahNLgUaFSHhZmzceFvZIW0xIbCvfxbRr
ttPOhpyWskDN6EO2VtGXHpami8WshDM+QnyQIJhntJBk8JyfIHY16moD8vtzzQoQpVJKC7PM1pTKi92A71kjO+8nEtdc6uQLVVZSZTOQZ16yR/2TbTI6Drvq+4g8mlDN
Dx1Fubaiby0lD3gxNOL+8mq0biQpIxSt9ZXY83dP/7MWMqwMTSoXUgedLRHynAiaZWFy//IrGo/ElY1vBzgmf21N3s4fgHuMGh9mgs8Hvwgi1OF06J7rhLX/L+DJ6Wkq
wjRVVk0xRO39QPCCXzEtm2pHwe9FvM4tZ0+MALM+i6CayWn/1EJx2Em2c938CLfdumT4kmJUVhMG2UlWgs8F4Bv1NEkMHf1jvoaoAC11nkDqUXSTZMTboMxo6UUD0oEy
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereV5RvcEF36xphpld4lpxrrQ5f4n9Peq5G/nDUiU5kUNUE42Fmdxuoj4WbdAfPX4gI
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereV5RvcEF36xphpld4lpxrrUhNfcUhk51uDnhGxcZYdkM1HbniD8D4bqdeoA9TVcHc
9Rl5F8a4M5w4pRYWHuYaUPy5ytTi59N7FtUxqh1dDgTBArxfC3ge2ZP6OrHdyfIs7ycS11zq5AtVVlJlM5BnXnMQFIHq5HkJID18sbqS6SXpKkwaRiliJTWsb7wjD0e5
v+dflYKzwLGqk62dtqauGyzsXxJFUKc6jdF8l32cq5AStlxy/p4+6JLQkF32FoZFeQEy7UR8erpWbbj0KjH9x/L/X4mNM3MqcgjUVuuK4u/+2NEjqFLekXbVejGoH+gA
mslp/9RCcdhJtnPd/Ai33V3t6kd0i+VOs8txXR/H4yAlDxrWsyXMAHRZcgZOzAl0OiIYTUpMQTLytyCCcYUyJFqgBAW346l9gFkARCraKBscPYxgbcsrr5jxZlBdoDjK
W3XESP99qbAM7rsLxvN0zPlUdaiTHGfdlupxCz9uAivBArxfC3ge2ZP6OrHdyfIs7ycS11zq5AtVVlJlM5BnXp0MaiaWUSAZBxVdvM7/R3CsrEvqI+xz6jtYNjO1LoPs
gIHIFUDkH4IoQ+GgDr1NGT5+/uStayjc0uWse0YEnwZ5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t7jn5SxzdI96hYBnKV/WP1e
NyUT8rnVO4rUaPkun8OIvH1rJX1Vei5lbswrpmr109h5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t6JuqOihxHiG/YzL1Yb0NKV
p8M3UrFivGVVTVns4Jd/is67Sq26hh4ygZrpxla9/GMsi2fUI85iFjNOaW1OnYnTmEEWfQxbP93K9ZXzNLiZehXJxE4DsGQE+ZpMTWs7qWYztNWvLWHiOw8e6KQYqiVV
FkmlRKby4EsMTParB1+N6ZzKnEXS1DcaelQAgVYLym1+TGTSSYiAf6TiBq5jwH+z5+/BK8A/RbG64eMqEJu0unjoGVW8T2R2+6QowZkYtknTXVmguuTKYmWBi4iH48KW
ksMqSiifgqtTb2eUoBoOFBonbMo/hCM6liIoK/TumSoBsYi80wujwYmZOUqIX6lC3G26olcOfJccl4+XBcSTcj+1JXQ05Wp1sVCexMCULSIdfdvwG7zENHY4pIXCXV2P
UezMiS+Mys7W3aT2xjIbABrlBDiScTx5hBjhMWL5pckb6nF01SopCX16TCndYmHX0cFCAzNNXKDi448SDuq00bur30yqmeDrn14GnYPXF98rZYCUTFYMwF1wG99nW42n
gVc4PWPtONU6NSARoPa/RadHsyoxwuFV3mrbK/C5yEl57kBwWyUnQskbR1h3C5GWJ+JXuap1RCxGNJKtC3g0I5H65hR7gGHM1gMeKVASmhhpxK0UeZmhxTwABie5qd5R
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere3F/s49eyKZoUk/QKVE23yrsbR+hOptkb7Sf+7T6tucnqyjzqbEZbb7dxi/H6HkJ6
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereCnOKA91yt1CW5nUz/lGI3aTnabNxb2xrs9BhnxVrAZpI9E0uezpYuQcM4i/JZcwJ
B9qb5n8zHUqE/6jogl3NZt/0nUy4+QG7Fh3B+DLkzzCN5pgOi0f4Mhg4p7qZWeJC2Rrm2ZNv8+2f08URrwfIDZXcmbAZ4CmJzFYRFji7pJEgTlG3/j+WSqBfeTKh46y4
spAK2LA7QjC7Mi701Fjt7noV7uAetZlJOdVtHxPJEdaqAsro39fEANL3gGPr0tqGP4vBXWptvaQglP9Im/zVtld0+YcxGSNw+8jmpDma0p95/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5U9I5MylpWPOOXSryStIt5r7mR2phB3SN8raL8rU01HxGAORuk1tK4mlPPS5ODjtJ5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t7uAtrr+0wOzzJQVYP5j8y9Td6dVkgDZ4ARz4f6FkmzXY4l/TbIU+DWxXNxC+dKUz5YUIca9TByX9BM1jvZoaUx
40p6M+8SU8PJaiNdKAM+RUJu1zqxD5DPLm4ixQRYfKkTW8h5u4qIrb7BsQC+T3SHP0FDzYpiZRa9Or0LJ47UFtvaD8YuGYtdyo6tJ6jeuQL0FlG4XRrdiT1+SPRQTyTY
8lMt8iXpkb7L7AYS9610/ENGk7xXrl1XlEdxfghD72CHlqQDZ5iG3b1SUt5AFotKXD14+uDOwrOt1mpJo2iIyl2rxSyR6dRTi3lsVmcleTDTQJXbrgqO04YatX5OEsos
+AXVjbHDCvLY/XyO8ZA7U62Q1PJ3dn6l70Plsk8/EZL7SPIElaG8eKtARzhE758ysA2FvBLFWcNh9irc8XajUynbVeXcj+J1VShYS5gdgY8iKI/WfLmYRhybcmJZqofM
knq3b1W+GzzWtjFBNyLl+KkXPcrYhXkrwWyDXT07jo5+2dV3XkAPUJkXDa0vF1L6XUDqKyVKR7I9C/gVL5nKqI/ylW6ZargGO3m41FrMdTIatW2/+x6j4+4Wq129ww35
qHYKo/NjxEe9u+M1QR5F6OJ8IffpLUmhjEnU0XosPECbhZTTj/xkU3FZN87NWGF76BQSfXJtcDamKy9PIHKE1Udfz1gmESYe20ns8WoX1/NKqI6+XiWgALzrfTBkE/eJ
+4R3SJdSlKa8UJaUTWDA+nm9Lck8WoMumBv0m/OY8J5bwo0KeuxVzfCMbSnm2V/xG6m4sIyJzdZL71k3ijcTDyHEc1lPmJlCWJ+aR7QTxUprQfRyK/Mt6nmcUv4oJpgj
B+v6SiOMUn9UagN4WiolqZ8rSM7OrDIJWgnJYHTyuasVhVet98W5t23ClKPl4rclt40u0HgsLNv4TtFESi/Yq5FXb0r6fhtIAuNvptEsK+QZyyDvYypTTJKHhJy//1MP
FOftl7EhiqX+dE8NHoGwAxErSlzE2lcRyOdn7ra5HBtfNA3xz39PtELFVRKNDAPa3gxXdyaYZyQuqANaZtL4fNtt7X713eaq3AH7Wqj5/9ZjCngyWMiP9XBuQt7/GxME
5qQEtG9kmJLPQBiYH/y3ZB3jzRbGE83iZmbvM9MG7UdzeIkJk8cEv7FQ4y4yMsafOmKIGj99FJRnC0stg77Q5saWlQSVQxjAtFXMYzIh4IWYWy3HZpVJpcbQDNaFQK04
3O7L5gQ2pwDMoqUvQOF7IMAnKFvJhzL2o0uXPGElOLoEXlIhtQ9U1HLsHk4zeIxA/5lEDrTkNpzc1m5L7t0ghgUfE3FmUfY8Y4vUJOjd+XnJvZ63SZPhmBKALcazPoLv
ii8MvNaaq4RVDwJ2D6iapYUTjW0e0gobr1oVkxdg9wfL7JIvVnN2YTpenbOlx7hVBr/Zj1HIMoS90bdjc8iXxn5od0FKfb0KTnC2Y2KA4vFzBFpJvxCOzpqTPv7XOYmu
D2Ad6rwLd1J8zbiN8qBrXfjqDiqSwcjXGI1KZY8hNtZRktCoCh9Y5IhCfOoOwMz2fcPd8T6imXdks33j956TehErl9b5kzHzlDk4TyTeYtK/faG9z96lx8ObkF339DG5
ML1TbCioXzPqQHk4NxH68vKunMRWsaLkELmDyRwItTg+JXmIwuFboBO0KDDHhP4e/oGziBPmsXuXoMVp9VnoyXO4GcYJJY/G4Zndi780nRE+JXmIwuFboBO0KDDHhP4e
xmpDqYVkKN3zju3ui0lTC7DZC5Ppr/IyG1TPkf8F5AA4fyRZ/K6RgSWnwHrgbSL0lUFlD9ytdWEW1SHZ/Gl4WnQ/q8f4/ElkvW/sFUvfkAYLeRFLZ7eKil/0T64grgcz
PzHJp8jWZ/TsxTv+jhSrK1j0G/nfAg/QrFlszMkf9lf+K43+doD6MFW45wjbRTyvgmIQol4ARYayM1HR+Rt+yX6vI0xmMacLvrxvgBTipRsdCJC8NvZqLKv3mXT0wFV2
6Z1p+rySXueGzTk0XSPwwjOiHyOnm/u0S95orVPQ4lfUnkF7A5ODKb+Cw+TOs3XYKGdEY0qhnbytkt58Ph4T5Z20/rlJPJogScmn+eGEBcV40Gsx26IwW2u2hOVTU115
VS393O2Xb5/TdT9iJ9mgNbYWZ7PDTSsou/kaHPZ3J8EJHRhE0HzfCU1xb0L2o9Fd/0pJnA/fEBuF9YXKeeGyM98w0ScKQj6ug6u7NASHdgRLdEvQn5b7Lc6QjE/cYl93
vlLDxMT3jSi9P1AmPVD8hP+YXPS5zhJ/+86DUw1Ddz9pb2IAwPZj7Ur+T4UBAN2nDSBHoLQymkSEdbq4LqXjZaTXuw3dXB+zFAqyntqUTuy0B+quZdkvzVUdKdCpuBRT
kVuZDy2OuTn0fcbUU6v8faPjBLBY3Kka6NhTBwIopBTWNXlYtYOzl0zS1+6KjBkK+C4CuTl2ZsXV2jnJ1+eXKwq7AF7+aTNpghc9i4phSphDzreweSKSZXoAEamNvh9p
fbu95JYsKhBpoJIaW9M8ddfnMYApZDldg+kVu3dsshqYhhwpWqpOeZ9XxTiiJ8oxcXMF9qjGNmPGiKY3bGoQR4N4VBBsa8z+i/WZLN7BUQdPcEGaNRHoeQ3Fj8CtTjFQ
WtiJiSp6HuJnHGOASlOfzWm+gFwSg+36D0JrxHn0xkVMTt2YNbC0cMY/FL5Hqss1Cs7lCn3fau5D7jPcc2zGGerKPOpsRltvt3GL8foeQnp5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t6Lr8r2kow7UuFXqkdDQzjPHgtR5q1pjfdjG4l7qkwETerKPOpsRltvt3GL8foeQnp5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5hmgtklcio+Cuhhw3FZOS0tyz1EhCgE7zBWP3vSexc8c/MLYdn+WiUxdA1/IcEG+GsgMJlhdtacgkVHxNhjhl2
ZtLSe9x1Glq0D8kdkgxO6BTvx0jZUxafpIZB8qAc+VnMEsypj/QGI6Y4iUeYNGG2lxyoa63N78PVgga+PlF7vfQ5mVl28VUhOIeyVR9sd3V61YWi0YgBj79npBBMJhtl
HHu3N1PYOXJs+lnoW18f4lZvOINxziwc7tfVZYbaDNHJUfj0MXDTk6/SRvZb00omno0W2ggX8TKXKc2SS30bQL4ymsI5NXFCkbD/gE96Bs1ERuUDAR3K92b3IRXwamsI
2wbJD/oLToNcPFGymL5ELvZl2RbjSR6kGtcEOiXa9SCGuo9EAvAA2MW1Gkp8G7eLW3IlXP7P4EuyvW4zetY3W8WYLk/FrBh/FI6tkOCLBWqw2We/uMNcRJAKmeRHliCg
NEEJYerBu4P3objQ7RMSNwJLiRHecnXIe7fSTYQ5sS/vgx4jQmGOjwkLI1YURWWIlu+KfKJBjAt8Jsz1J324YkegbG/8B6/xjM10t6uQYyZr09yLUeKzGHpQ1sVQ/FTG
jLdLKlzAFnjKRjE/x3DTaxq9N/ZtLfEI+F1+g+WSIluTKRYJo7Ey/pjaPfDPwb+AtIoS0OOeLR+KHxW/EjXEsB+K5kVB+GebwdctVGTittmAE2gbw8eY8j/ufIF2z9Xe
BCPiTIKPfoVZzjuG9o36PPO0KpjJY53B6Y1WpK+ij2eFyI6kWbRJIpt5Shd9akRhumT4kmJUVhMG2UlWgs8F4HB12on+XPtOiK1aVsmMP12eGK+ubjDpHLynGKUKGwdf
aa7R6pT6w3TwWkvB3x/hrIaXKRaNmCUMeavMQtZW3HJX/yF687DgzlEKoCPZv5xyjLdLKlzAFnjKRjE/x3DTaxq9N/ZtLfEI+F1+g+WSIluTKRYJo7Ey/pjaPfDPwb+A
tIoS0OOeLR+KHxW/EjXEsB+K5kVB+GebwdctVGTittm6cLNhRxZjkD7Ki7EUsznhBCPiTIKPfoVZzjuG9o36PPO0KpjJY53B6Y1WpK+ij2fFPyIw8HVfWWN+QP+F4KQs
umT4kmJUVhMG2UlWgs8F4BzbH/b2BiJdep8xEhNlABieGK+ubjDpHLynGKUKGwdfURVqU0Rk8zoz2Ryn58eBSIaXKRaNmCUMeavMQtZW3HJcSavJQGr6Pcl/Q4sLhBcL
jLdLKlzAFnjKRjE/x3DTaxq9N/ZtLfEI+F1+g+WSIluTKRYJo7Ey/pjaPfDPwb+AtIoS0OOeLR+KHxW/EjXEsKNVO8X9+NFe+cHCE12P77+cExevyq/3mFRhEq4Kv3bB
gKa9Rz63AfDGH/eNcG8uVok8H48oMbWBX5z3e2stMrTl2616arDlYTtY6G9ujqdRbFe1QZ++wG+lzsNuC17pkhlm/vCqde07KV5gWsuV2VJ/NufjaXtetYCIPqLE+hlT
OtkjJTFF+1OOYTP6+NRaRLPpISpLtLjw3WISM09acE0XGjuOdvx3qok9Qvq5MBWAB4lfTMHZgnsiFce+ltqbNDeBfsd7MOgPbRu3f5qWxqQ/kBaElshPDg05+STjbMIm
P2yNTae7zI3+OYBHKtX5gT7bS0DF0oQ/LQZVDsQdWjojs1gU431w+g9fvSXMwq1AI7NYFON9cPoPX70lzMKtQBgZX6efd3vIYcTz596weGk62SMlMUX7U45hM/r41FpE
U8U9Gdgsl2bCCyNt+jH4zh/uV7h0RJGy69huyCm7FbHL32GBRdSx1O/mp5KnMvmSsZfTHfsR6FSqlIcLa9KzLY9nrXSStfbO4xLIVN0d8qE4LAwWmKSbFZZYwKqSMnyJ
Gp6BACZGSbg8E6JIMXHvB1+BbS+sxjA0uypoNEeHrlvx2CfuSuWsDwPezw0gcb3LUiuQw1HiHElcHQO0009QMLRHZ2OFQFb119YgzhrFjvdZY/GtuYd0FXqMaaGXGI+8
G6suujuXVufWlqF6fF8OPeunrLlskUmBlmGScAbQRULoPLl6j0Pg/s39ljsaDYPgZkMWVrSDimJV8jPFFR9w5T6NUkjqkMkkMdIkBpqEIFc/kBaElshPDg05+STjbMIm
nBxrz481nHfUo9G1B4iYeISwUNsYcTLDDt5ZW7KCRd+82Frpb0QmXJzZX/+mw0O1B70u8ulMNa4zvH0TdwO2rA7BiHLPNTqvgYWYjdBg0XZANiDGn7JIfCZ7GmtyhQxD
OhuXG7nQPSHfQ0Vk4AjJk+ZLH3HWFHdTfICOg65+WgOZ/UQKjaP29R6XNIKp0uvKXRB9Q4zbPYCUng75Feob/l+BbS+sxjA0uypoNEeHrltfgW0vrMYwNLsqaDRHh65b
8dgn7krlrA8D3s8NIHG9yw4bCtz6HVsCDnuM+zs0fF9jtDezIy3JvN5XVpkSIkFIb2Qs9NjnzAkXyqLugCm4gRBIbQXkoDa3pZ5KUvIMwYyM3W7Gqpi1jGTASjaRS0UK
ZkMWVrSDimJV8jPFFR9w5YlPk+jZokn/UT5YCef0qe6mJCKVNl3PfH7OQD4IAaiYbvxmg4z3m1NJzR//VgB16dZeUbDgj9wuelaFeQUa63uLETXLpLonrtHNaPDDAUic
RmDRM3lw+BjAQ/gh5lH8DtJOVpm2+fkqzqMjojydTVlVEkw2oznH2QFAXNPJUNTu6D2sc/nY7JCqIFA9/NUGBWihqhLmDoDe06Utz3dUO4kQSG0F5KA2t6WeSlLyDMGM
jzjsEXmqVvpx62dGJrnNDFCc1FsWxApSkoTiDZQ9poSlWPQNO1f45e0rVYC7fNeOTsL9QI5xodUQ2tsHm163DLkb2Kmk4jbzRYHhzu/1Hn6mSxk36mwWfOcywTg5OpXf
Ko4WgfkmKIxoltqEn/XKeOg9rHP52OyQqiBQPfzVBgVIRCW64d70e2cpTHKYVgL1PgVQLrTRy9hOSEZPuZo+kosOC4qcuPt1xK35cTunE/B7yJTm1TnZnUAR2A3sXJGa
E0EkkBFKThJhjy3RR9kCXURG5QMBHcr3ZvchFfBqawjbBskP+gtOg1w8UbKYvkQu9mXZFuNJHqQa1wQ6Jdr1IIa6j0QC8ADYxbUaSnwbt4v6hx4j0QkLS8PLiVGl6MMH
it3H2Pon7SyzFvG5Pqmv6Cb6yCcl0ngrddQ5azFTVlnXuLbzulk5jRV6spYvGDzbIdvcdnZLKI6dV29qrVvQ8qiJiswDZE4MzkuPA3XFil6faSjTB1wYbmU3eTTHZSzP
s1Zg+naVG2BdWAPYIp7kz19uVKw3g16KK1fZNNrUeJRAoxbrzDwhXccN7wSeM4p18i2AOBIIf/pc1rZImbk5UyoaPHzoKswnhOkAZvMVMFuB+vpO+cZVbyN/yStpIdc8
+jP629ou1aaLHj5H0wX+Le8xfhmtwhim1vRv5Gm/Rg0miUWV3hg0QEtdJhp2KP5papdkUSn2Zc3E4tIldUvZduCIr5oQUhZZolc1w0s1P40qFAJYOBgaRBR1aORvTiZo
eOvAgQY1Vmvol295nhhnH4zvhNBjom3yof/C/VKAUwnGAg7aj1+MesywA5LMgwodChHbzwEAUofZssiWPY21Mm2ZXpYiPEXIIb0uNgOBMo1Ld7Om0ocVEwf7zzVEpJSr
3pmaAjVh9abmxTnHuysIFYH6+k75xlVvI3/JK2kh1zxVEJnuP7c8TTkQn4ZHpJvAgHHkVkqo2L1z51SCKvewVWJwdMUWq09DBUUHfH4cXmW9+zcwpGmFZxG35Ri99DP9
G0U6Jfsz0sUr7BqPDxodNfPS566q3j7/wtbBheHxi5x9b3iODC2x0T0utsygw7bPuUrnFCB66TGBT+UXv07LNkagiPiHne46oJFafv4pb1NkDbLuelUhmZmXhCzbIK+S
HKqJZG3Y7rLMVq28R7r2uu4qDyF3O3gsB+OsB2HuM3tf7djTBUK6FA9Y2k1/4MotOdjGYv9QZbsbhMROBfrZaLaxlxBzdimi32cdjY6BFhlFusaL1ZqqWktLzXW0kgbL
x0QrKT3qU16bl3EKsDuzsT12F5wZQ9OpBRH97dSJwCwCQSmiNPwATbwOLp9NVXzb/eAEmtSIRyc43KiNiCPyvmOyGBzliNQaihNMEP1+NczKos7TM/Yk6o3igUhfrmDP
CQMkXp/6uOx0DhV+M+VXgdZUH6LP/ieB0zKjf6IOQi/meGhfomXATHVN9mmm+qrlDomt/JmUrroT9CtIuYJPQgbhswdWLFle7cGDm1c3S1z16XWtxu5N023G9WfOcRaC
+3r0UVA6Bdz51Zmk8AMiOEsku6m5koT6b8g7lmaTxA8jjIitqoQJfq7PuoNjt/8HUNJt5rPC3BW07XYn5JvJ8ktpHyvsmOS68u2cHjrLDKVRmTufiQQZV5NnVYegAi4p
dbfA9s75fBbFxqyLLtK+22uYhY/VCAbepYxd8OXXugd3oJdd3aOvPynEYmCC4Prs73+8k0QPX+nlc3lzbm9aUNPdYxFW2xb1tSUA6s1yW3T78YmN0Itloj4Vkuh8GQSA
tjxEykUv95RuZm74PMyNDMuLs+wgfugTm1VXgK7r8oC49k3RgUXemjWFjdJS9kTYl0T3cVrWf1DEcoGu22Wfyvnkb4O+a87BSoq82rvdhPWqPpDVWqVVsclJg1KYpRSb
gHWYV1tpk58R+39FHVm3dzoy1SdDUPIR1bKkC+ZDaIqCv+MvwxxLYa7aOm0QAGEE8fqHyYcpLPUHkkx5i2RulZ4rwkhxZt7u3QCoRnctu6e74wV/ZlABJu+8GJc7gwQ4
W+wy18PpbfNzCBCGFxhLfJHnl5ZpAZV2BTEQZkyQdQRiAvCwRlbklYgqoC8x6aMG1N8rV6w+GesR+AXjoa5yO+8Ruiw/oCiieliU+8DN45VZHF6JVDeWeoKxTJfGOjuL
zAPd1tgjQPaXcRA89/Ycm1BfYTzIFPmDZ/z1FADkKYdRM8BHWmSmxh2e2wQmbUD1JJpeiwjqjDHcfQAY4RSyFMZLPg8Eea8RAtN6dn8fhHEjVF1olgHhTx8PSsiTYxgd
TGEyRGeslm/oiuevcE/2y0LI/c5jOkCoBx3RNkyo3VO1QnHSKscMFTkuta6BfujARN5jwAZ0zk2yJmJtNwvFVVDob9NPD7OEkIqnVGTc9/n9r3X4iUp4dvkw/kDTSPNK
Hqk+JizfbYE9oFkYjsBrIJyhA0MMehqd8n7gDTimLoPuhCMDj8KRHIqtxSWjAziOEeD+NhmNrnJt1P91MeknIxaqZJFlHHL1D7kp3lfy/DQQhWnQr8gzLLdxHbudR0G+
eWeqxpUEhVTHXi2uBN240OJKkOSfnUa1F2J4UecceAb3CClpEpczSCjJ2oCGMRIgl1oyyVdTr00hl8il+5UkV/MZ0hGWudOMP76eIdTbMqFCL7rWl+P2TXDcnzKmJr0B
W1s2xawRa9FU4f1Wg0+xvut4KDH8dGudu+AQTVTnSopwxsJegyfn9PIF88dceJoYzqkeKsc/Tqgl6QoEjEW7PqcgSH9rwMnsEd8/Zh9D7HaePTTPgSBrhApeZEkjUSZH
WL8sooPCwlKdiWCA4Dp+fMTFLALMBxTd8Ke1h6yywattT2biqUD5+3fVMYvi+hbHvEKlFeoKPmeTuIHtLS3TlRcJwhJmF7BUgyhTsMAwqrAHh6POrpkMmHqOurR4BT1Q
yzg9ihu1oBKf+/yui4vPdO4wlup9jCiMF3Sx9H6o7gwj6U00Y8lDSIWHZ0/9D/6jef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ilQPzHL0IN3joY3jfA0luyqWiBYrIPb2I8ceHZju1ThlsMrDLiCSCoK1YpjfwRWsef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ZSfJdJBYrDoLZ16UTLz3AstoaG2bnzljJCqOHh+Ufxo3CdYY1mHbsZTBljfAO5/KUItTN9MlTQwcZDn0FqlMjypr6V2EaUyndVtGnHTuIeAChDzxyU8+YTSJbJ/ZxRLy
rwsqt4ga5dHP4K5c4lw6+lVTpHrt7kM0L+KvIrFl6XBK/7nTIe+0iT4Fvasjt8OQKnWOx84VfMFpRkXjyZiO6QsZn5y7s1VsW21SUuAknG8KDLCp2wOrgKyNDQ11aVp2
lDCTMxU/qI2Rlsviv7D2zDBMpSdx9Cpg5nZeB10xv1gsn+2ach4KHRDRCyRamSdDaO1ZEIh/bEY7cCjyrR8jkpmjTtm4WkYOabp/VW4py2o8G98JYxJcxQotSojX4fiC
lJSZ7sYQ132QUjB6CH9f0PuX+at4azpdVlWn5rbcT9JUN5xcV/20YAk38KC19De+x88DLRoMiljb7JEKYdv8QVN8bQdxur4MfDo0FE608Zu86Qj85pgmu9LJdf9d6p6z
sOkIPprIv+6k5yu5q5FVOLoU2XsxfAULX+53qYzPuFZsbR97IvAr6rZuZhiPBUnr8Ooky+K5/uiJgEWY9676ThWqPxIw0dRyvpC+fSmWCcG479twGQgcfguof3RXHfbU
xVjQlUVKKDWlJMhudXLm+2Vwm4QOup/FGA1sP/4Z9VoOrXxonAPuDVPUFLI6OQZAlQ1V4tA+tSVAYhkymIBTGtS739IwRBzFNetvDGgvGXKDjNFB2vhCmBvgrGK3Y8jB
Fs5thffydKelMnOm4do64IPfqKYZC3Tve5v7rPSLGYGlsfNH3D5TPSNmtw8BrCl4e/SeBYHW2jU3cus7VAdOYxBkEqklEK9TMMxV0ihzHmakQKrlIHaBI9yZ3L2nkeJX
Zxba7uuOgJ5xy/yaTYw6dAoCwoGLus5X7/d1H5v/0QIxF0wU7W0DLDSXwB9Y2EqJ5WJqzBoX33czvvVakAOKJnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3leUb3BBd+saYaZXeJaca631LsnK+bfdZq2hZ/iiZvef5ByVkO+ApcDdhs9rPSu0TiOn2Nw32BeZaOwUqp7Yp8J5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t4y+MPeZAA0mJ2FXwAbXovoqNIvWjUex4+ce7/fpbVsy3PSCnDq+RmclDW3/Q8yc53OyGD/3mJZX4r5IebRCP+v
MF3GiN7ga9fNaCE2BnGUXl1M1VUrwiMkjeIghg8o1yhrMhr+uOkfRPAadFFNiBSNC3tOKoQ8/o2hAPKYHaCRhaJdEN0gOkhXcB2bJ/KLjQ/liXpEUQj+Fqep8og/06yG
G1eg0c6QzyBhiBwU5Kiz50i4Dz0Bl+Wwkhdde8G60cokMZqa1ExFTr0OowbB++wTRenKeQQ5RRYQ7P+l3f2ZPV6JG+dT7WbZdcuoOOUFXOdI8ovjfh6DXMwCZZAjjs3m
ltr22Q1Nfci1zgmBOhD3+bmeOgaMFQb+d3zCHlcdaxG74wV/ZlABJu+8GJc7gwQ4Yk9baK1R95RzEsTIWk5K+kR8L23PkDo7pTAZOwHq0SFPHpqwBQNJLqanqrrtW0ZU
vjfnITCsHrfhMtxOduFURELE71jrWiUhS/3lpsm6n0N3ssJLQJofu5lLxiXqNmPAmBE0dh7avYN5M33RgcM7Ad0N8JdZ/fJAiZ/OevEQxsLZeVpUEtML/fGLt389ydx9
j2PnjKkrkTwemlnyLsJAaFhvKTmTvG2K1ogy3F9sLX5gviVlbnJIHk2EVa1DfA9KuO/4fCxWfgw8Xuc6OAyArTen4HQkYpOKo5nPR8R1lsPjZoAE5cnd5ILQ0VjQ9vpA
kykWCaOxMv6Y2j3wz8G/gMOG2xGt3Vhu+u+WykYo9brDNo0TEEzCu0TK6oOO4LaajODGvAk60WkEA9Z0n9L+zr38mxw3oTDQLEEtvgGxNw1k06MmBwmRU4L2p89QEtyC
BncRGI3irqEIAyIDWXjhca/L41rQazFC3WykIrvLWFEGGo1aBbtfYZGEdvg9w0CppWgZd7EZ3MRaJzgh35y2kDnwwKEzePot+2TT+uvVw9LK6zAfSh+dtFLe2CB+eKup
XshRA6fLSpTK41oG+hNAc2thb1+a+q8sb2amdawswQ1GxIPo8iU7ED24LF6zKq9l8qnYXbJrqOi0st/z6a6NvcE9itQYNqc+yJkKK/JnLm6jM5HUZx88urGDNVQPA4eh
vETXqlv8v/M/HxM3K6ssVHpJO248hNvmGW5qQMbZAsdOgwLge0Ig8xjuojgktEW3PQiELy9rEXKw7AO8uG7FvzVzpq7S9ZMY9lydATKbhZDGrHicKND3tNJZNaDRXTMR
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere9t+VOOwg2pHWjAe/PJz7a/rO3ETMgpYNN9QFfFk4437MdgSprKG9RL1101wpJqtS
oq4kBeMStmcs1OuZ1tzG5K2HygTOPRXllHjp5s8DRHXPBuYAWKxr9+sMpCzNrGMeR1l+zpQTB1ipSsx5HD21wKCy0r16TtLhCohBAwomqCE1Om7RxjlppUKTpdPPSuE4
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereFWRD6byeeowGyjZGbVOjA5akJHmytQWwHaCnJRrCuC2pGHKGbhcLzzcJgqef5+xT
QjfBNDGlfb07TH+8zkcvA75n8EyR27jE/FwxZrsI+NY95Vx/wJPtNtofirkSdlMUGuUEOJJxPHmEGOExYvmlyR2GV2bJ5VwkvlYocyW30LGwDn6Zqk1sbXEL4Dl4GItE
QnSONHGwG7iClx5XRDD1bfyriNFrWnO0BX960XjLK9ti+NNBC6+bEkEDubXS8qy/o6Vbkr95+LQXk55QbQ8Lw58f7fKzwD64uHOuwR+4wDMUzdKL4tlTT0U4tnHWfWdL
kzM2cw6F9BbfX0KI9FJOFQZpsc5VbUvgLoP7Zz4sFPBUgHo5FkyB3G7t+sHoZYHeXZOmpJ4X9msFwXnckX0liKGnsBlNouNOrCLT2P+PANL+dodX9CLxGB+SSA+/IudY
htu2ClTTYP5cdb1g+U+0gZgJlMcE6uoXHuZTDrtIkbdljVwOMM6/GEpI1cA7GCCYt+SsEzJPf3rdxkAPodM+akrIpsDa09TebAIfmOjRKbLRwUIDM01coOLjjxIO6rTR
e5SJk0if1rP9rswjpT5TXNDesVS2D8e2ojgDvnphFpkJqy1PJvdHFs23+0xPW+8R0N6xVLYPx7aiOAO+emEWmQ77I49Ro1GfhHryFSmIqtkBZ9yqnJPk5r2iHId/kab4
WfT7nav9uw+tgvxBLdEhg3n964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3q2xzG0TN7ef+5Vq36xqt2CH0h549QMnl2W+mG/uCRC9
hdtAy2fs5WDzQg7ra+63cD09fnmjPkzjGI55J2cSwfFGuae4fGEwenoiYdaFikxtdaxhM6lXP+GrcfgotMGbeve7CyYfSjNXj+q3K72eAnUrhG+58ICvDhf1olB/T8on
Dm0CB4OAGsbMJOfv1npeMXn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3o35a01tqRpuz56rLtSbM6c85UHXkPqMMwAS29AuVqlz
FUVsA1S4QmKDs0YXBMkOGw3DzGohwlH/ftsFOSCh/kNtmV6WIjxFyCG9LjYDgTKNRYuDkCFM/rUnmS5Iqs6KgUxjGv7138coJ+wAoOeQB8IkimXCFZr4lO6lo8LiEwBe
tw+ORuKuy+MrcMyNmTX4BZ3sJm1tkCCQekfJwMJ+JdmjDoF0imH6Tj8gdwGRT3rVTGMa/vXfxygn7ACg55AHwi5eqVzc8qKRzt1VOHULYA72jBpcSnrbxD4EVRgUIGef
flcQ4mnFwV+eVN/ia7OsjYxxIbVbjTYsv7xAUx9rTU4NIEegtDKaRIR1urgupeNldHQVY/Uh2nFjf102PuWuOF4vT4eZsCDwypIzO30K0RSwMNKbaxid+8DHjspBv3M9
N4KnMtH58zY3xGwjDATxbikrqPYJf+ADS96qTdpCuDFgAB+AMEsKyPQo1MAUJ/RKOI99FZvw0YJtWQvFbVCb8ShSHToAOM5/83UbHO6VvkfoLH+c7kag99aCMcsft5AX
iWGkdEpVOHnpKtRxDXcBw2gT1b8/7jLpW5tdS4XdrgLAvvR6U+MDi7IEg8YgX163PMEKKRZVISxsxiVf9uMsoOdHuPHFlruBpt9SrrPFFJzk0DOnzEH4UjhiZYRmlpkW
0vyRk1PzLwylnFBabBQvbgEM7K555kzAavgtPzE3NOpl9Z/h5jaXsagWh75/8Qne509k5vcFEip6BhvUN3UvUrwI4E+LehOX5cHuXMHC04fSv4f4e/QF/nJ6TG+RmK0q
7LOC2RbCc/4ZKKHs7iQ67ke4mBMy4m2Qp4uf2JX5gDRf7djTBUK6FA9Y2k1/4MotAWTZQK3OZVoI880U4UqGqV2TpqSeF/ZrBcF53JF9JYihp7AZTaLjTqwi09j/jwDS
/naHV/Qi8RgfkkgPvyLnWHz+u8Z+jkhdL2aTBD9Fom20LVxTizXi6ekYhDJWBuryS+eKKGoHy69+yi8NRd3e9xkypKOuoVOQsq/r7lqDuzOFZXi6hkxL+5Q+0l4mAJ7G
/pT5d9Ybxqw1amDXHQ/9QZ4zXg1K/ud9idWOuuonZRePx8v6eS5q/d+JuVeKT50ywVwkpWADQw6nkaZxLfB47LWyAElAccj8u1cXM9nkpaBq5KfxNfeo1hIpJCS/kmNR
sxZ01yTdd5hbmTr/ie47LgPUqDW5ukFAnwfTsTEc8UUinM0j6wZtVpb2bTgX5fyupuJAzV3naFPk/CGIPs4NnnY0+yMTR6q3+UxfY5vPl4u6aSL07F9wqwc/3Dv47mHe
iiMpWcIzP2plnaQEvk25NR8/rfTdJMPxVR0K/sqxmpkruWvfV6jMUwFSSksDAG1FmJt2bX5mKTwqdZ3Kl7rUp46SNbuPQMqWtuX4tWsMHigaXroaLAjpOJrVbPNnKHOP
mumQA7L95ynuEPXUijPAk8AAzroqA+NDxjFQ+O2Wcw6cfQqEc4XBAtwxlnqoCgMYedTfzovVjlA8f/aPJx7N2hVikNDOFnQCvnLs0gxCSOUd/ozKJu8VUkpV+lnFu8FH
nrX+tUJ9xP62P0tG84UMrQFk2UCtzmVaCPPNFOFKhqldk6aknhf2awXBedyRfSWIoaewGU2i406sItPY/48A0v52h1f0IvEYH5JID78i51hj2aS6MM7dA44wKjqf5Ij0
pK8cyk8L8JsCO4D3KRI2ECMWQ0JSJvHIwupMb73lq+u/XChX+b/zaJtme1wSN8bEw4iOP9AeWOiwJUERin/z+siG0ynLuLFtU/W5RFd5FSoVA7kkUe3izDysyxJWvZ18
wxeeO6l3osNlpxh6Wjuk1WuQF97x8ZczvEM3kN9Np/M22hLYHOymCVriBxC7xVtHO3ViuILwqu5urDwuiGVoOwBXJsIRgCGyHpalVX5LMCFMyIOBp+N2eJvFZFi8euvd
RxZ7Hp1BzRW29VyZwZn43H6/+iWHPH8ntbemT60fQ7Vw4er3dhRX13xu591hpW3B91EHni1y4anfpy/dPmiNwac5J1LdQwzcaMIpSTxjgm3j3AVY7IzAF0oie8kd4B3r
gU0t4SJOrqYs06Dl4NeXiy53nN5tDgsHlvHJICJ5os/QJ1KCzdLouifr1P2+XtV32G5lNyjMSOMU6ezUHP/cXCIL1mUNpcPsjNDFUuD/PJ2Z3ABnmdb0hZfb5tV4yVwi
Ck0KqchT7iaNAKi5pRBpbmCisoIHCtr5F/NCZcbkZBVfiGePRu37cw8+P/9AK0qJXHa01zdbL+GRKa7srYzqRvDw/axsUBwy0bmtNxAKNSQfMvc+Qdry1iDdPN9Ym/Ae
J6s7xJQa4xkTUi2kD8iXrzEV6/qgYGZRcDFtChGgj37xwatWHUrvs0X5ius13YzNI4+1jIgfxLT2hQM0ftyGopPKXZE66yg/WZfPeK7mjQhzmgwfFErJK2HZ2lbWz5Z8
wlYWmNMlG7wg9ac0LlABYomsOHFn+3gpRdWpGUlsJzOWoJHv3AuGsbZ14DofIHYCW5YsvQ1AhTJSEqKsU8MGT/H6h8mHKSz1B5JMeYtkbpXis/zC75IC4Ur17hBdy17i
h0lrzejfrZsHdfTDfXtWDUpZCSguyF48pMW9E3qcWBPSYdgiIfmujZE9TTnge87K0CGJXNdDvMO2gr3tbqO5qeCIr5oQUhZZolc1w0s1P41yFV1Zyr0mQKEft5vVprGe
/fxViLQT5kY0NsWBXeHgVTuCG5c8ajvOYK0B7osNeHn/zNN4JhKKYnEnZOYK084GztMdrxWC6B+5LqsEOmvFDoq5Vx40PDp2KRHShmhDLfeqhjF4f8vbUPuTaRpXnE7G
nd9EVX9f4E1k8VgdOFigF0bw7B2IJl/04IGITK/hmMUsP4ScNvvMGfAc8aH1C9COx/ao43dVbsfBRtyk1COmZnRQ2Zlm0rzPfrTE9aKZzbQ+tGPBrsQVUsbYEzQbPx5q
2SxBVyI//OVZlHLGSsfrHnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3mcYtWh0qJ7wYPBs6+i+KSqemmnibnIbJcv33sKxYFFB
XdzEdSVh36VbCGg4iBzTJUJWADOoQavr+Gl0KvHZ4GxjQZBbCAaKh4mYV+y9Ly+Jef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
+UyFk/pXWElHAXEColod7BoX5vzI76+S0S5DF6emXZG2sZcQc3Ypot9nHY2OgRYZ8C/5rxoUMfqwRDk1U5wo0ebxiDhl9xKKpfT2N4NOx9K41ZU+z9CuZ+4oJQ0Z8asp
5PFTIrePJTiwpWw1Q2mQiDj0M3HnqxgVcXLVSCI0TAK6paskUdQfPKmu/Mwi9s1oWhECH5HrB6B4dgD7ckv+jWY9UkYRo5JjmjaU3W7fdA+H+bI2u7TkjtNIqR7TErS9
p5v4Eh4IHIMqkIxD5SnQrxU9LlbYmw+iWb67ukwiunTnBa663eZL+LhIMvJzseMtakYQl0Zob4C/D4R34pVrcsnSiUURZRXXNoGxHi5Du+u2L8NROgbDPmK6G7Cjn9Hm
zT9GefxFW1GF+YF+022hQ9sGyQ/6C06DXDxRspi+RC50ZgSHS4KQn0aEA8/4AGI+N2L+NNOcuJ+IfhzfqRHvuv+5Aj5Weq5S+Dj62m+TvBHk8VMit48lOLClbDVDaZCI
k2hdgjXb74PTysFoDKb0SLlasCSCkuctwk8iqXMrCH4A3csfigseBn8XBFYNbjGoTghOS9Sz74gH2McY169jJ0J0jjRxsBu4gpceV0Qw9W12muXavcLgawI80j07eC3o
9xNcmsoV1d5rYpGd7atttl7mR4wp+C+M1hsVH6cLhekZLA1E7JItKL4WnQ2ehoudgy+d+MAldUGvfzasI8Z4knPSCnDq+RmclDW3/Q8yc52MgUCzxsOaSFWGeNFoLiUf
pXc3R4nKMohkamQURszGNECrfqpV8sIZF9EDWGka1CuBmMTIhvlcI11ExMH501dZ4taa05zsFPth2Tr3lGQwwNPKFcReTMseGsaWU9IvwI1Aq36qVfLCGRfRA1hpGtQr
bTh5cSRR0d/DW33qqefrPzaR6bECs80bClEmN8MrmW97xmLLa40Pj8S8Zbd7MP6n08Lfv7kxbBDmz1rZOF0D1TzlQdeQ+owzABLb0C5WqXMVRWwDVLhCYoOzRhcEyQ4b
DcPMaiHCUf9+2wU5IKH+Q22ZXpYiPEXIIb0uNgOBMo3+b4sLoJMVFZK4J55CDFiNHQiQvDb2aiyr95l09MBVdh2GV2bJ5VwkvlYocyW30LGwDn6Zqk1sbXEL4Dl4GItE
QnSONHGwG7iClx5XRDD1bRBTB3aNGbZ5l8k4e0Iucp2w0D4bdPHY+rQGVAm0SpLEpb5QaX6Vqr9jkQ3XFXE9dy2rnpoHO0jHixvn3B+ytM0yuqskD2aEt3qxLBO1VsNq
o3nO/cNx/9m5eWZRk6FoxInSYOWxvgdqLrYCf9dGZ8cF3RiODTkLvfiqPH+mXdG/xdukSf92WddEvpNVSecFei5gUrTKr6zJ7OC11iho5HULmz4Oo2+89ie+laCRTX1S
LVtJs04yi2zXQXEP9HhJPhhNHCRoR5FGFKE8LfQK2CStsJp2x19fJs4WbVKDNFxC23iRia+wHOhCw2otFTI1K1/3b4SCJ+R6hHPSBztOWnEgyEUYYVdXUEtyhVhU//gE
kykWCaOxMv6Y2j3wz8G/gHQHqxbSe30ZjRxTeMgSQVGsUF57Dy4rLpUdCtnL+pLcvNvZUD8T03P9JU+5pde0NRCFtKjW1RE/nHOWbYtTHhZJt7A+TTIETPa1m2Dgn006
fo5hEVILghlrhgRzqQAbUNCfu21Zxy8KQoHZO+EFTcNjQCP1rsZN2fY8cDTIim9WFXflkGJqAvi16dtLhT+6TNfebF7abebA4EnY9xWCR3saF+b8yO+vktEuQxenpl2R
trGXEHN2KaLfZx2NjoEWGfAv+a8aFDH6sEQ5NVOcKNHm8Yg4ZfcSiqX09jeDTsfS8sD2CnH+VKRBJY+5+IcrPhqSJjR2XsOsWlezgkfl46Dio+dtFQB+kW9E6ktMqSuU
7/2jPsYr9/608P0jv5YUh+DY1EjIakEiWf2Rwq80oNad7CZtbZAgkHpHycDCfiXZ6TM6jdu5fZRZA1s2Cfbv8sHsA/3f0jkRT00U5v9ty19AUJoaZLuciFqtH7EJKdIO
JkQb/vWGl3+UWsbRaZRoNPmWUclXE6X3RILqkwTGSQ23a4bfmPR3HLHYce7W251/QKt+qlXywhkX0QNYaRrUK0xShCflN3d6fOeHSqoVRc6vFxofIEdkbzIidL6tVg50
CqeuVq85jBQibRz489/l5F4/HdKYCAAYN2nbG3abtSrNcr2BCFvCwfcTz1OaP1BAncFTJ5FoXv09zIinq0VEq+gsf5zuRqD31oIxyx+3kBeJYaR0SlU4eekq1HENdwHD
aBPVvz/uMulbm11Lhd2uAsC+9HpT4wOLsgSDxiBfXreavO10GvPPLMV3uJbG/HtwEZ51RUbdSMIIbJQVgw6B3iWKP8XCTLs923vdQGwGpGmzXH2TDiRGiP/kTlFYG5Sv
2fL8s9dXoDfklfelM5FSamY/0ltL1dMn/cWUJ1GtuB2IHgNGKgps2XPdShCMUiee68d7eRIOA7Y5tfGr9TUDy0QCcc029L4HNYdybhEL2Ss85UHXkPqMMwAS29AuVqlz
FUVsA1S4QmKDs0YXBMkOGw3DzGohwlH/ftsFOSCh/kNtmV6WIjxFyCG9LjYDgTKN/m+LC6CTFRWSuCeeQgxYjfKk1OxkkPPQ3OHWcJi49DO4IhnfEuhUnbuU/QVr9Nml
uDmA4ohSI6STd7GMExv7vJJiOpo/eC7oIe8hr0eH6CuJ0mDlsb4Hai62An/XRmfHvUz6hShrnxnC3E+IKuqUEv+YXPS5zhJ/+86DUw1Ddz+LlKMqxgR38gGN8hEOs+tG
PoI8AgU+qp9HkiLrUktSYmh2pbiRJQhQbdbGnFY4MPs7Gd/WQTva0+7HpY1MSZFg0oRizvhnEco9IqWtKECscJfMQhW3KV/qvYyvXfmAATQ9XIbXKuZoHlpnbeUrJA94
7v2y0qJ9wXWknm3NRBCVJyNJO6UnBLU5Fk1PftzbOClsmgCP7JOcj8E9o9upSZZaDSBHoLQymkSEdbq4LqXjZepB7zJV/MeBkhQAxuNi0ujJMWDeGCKggbOZN8nxX2gj
68d7eRIOA7Y5tfGr9TUDy1TPBNogvdszyvrJhJQFRNygIHu5iWbLq7QoIz76HWAQ821iSrYNVaxFOtpHUQuGUPci2LIhYe8YUtQGz6FgUf3Oc/RuzHLWvnK6SrHR5BKo
+bQ0UMB8n2KnVjI3TkdTI9r95nZBv8DTg4nxwYIlj2RfSvk/T1I7xU86ziyT13H2ZajnTM8sYfETMt97+GxG2NxFFYPMnKtq8l5b8lk5F/xuQ+tnZ8kpPXjqVsfl7AlI
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereYEfSAcQJRYoPsPUlyrDB5nM8yQqlDIQkTG0uPhoE3qk+dXNSfR0/65S1JaQ1RPkk
Vuyc2pAmAAAG/5D1Iwzzyr5WwajYQdrEZs3jCXB16T95/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5XlG9wQXfrGmGmV3iWnGut
UIpkKrROl3dL0leQiLrSlGPZbRgGZzXOuMI2ObeCXoB6rNRa0IvwvYT+SETOC6CElq8mXN+wQBp+ANU3upggFYIiG62QH0gX8w2EepyyCYstcqykieObo72dyXjtyP9E
wVyeNTQMiUfCm34VXKKgPyqOXw0m5vsYZf9ebt3EDEQPYB3qvAt3UnzNuI3yoGtdINTXgdLvEtTk+FdFBSpfl7xFOMHncIUa0J7BDwEnT022L8NROgbDPmK6G7Cjn9Hm
4+VvGe6rtYg1HmQQA1DsAvH6h8mHKSz1B5JMeYtkbpXkKNJuV3sss44CN4rMmf80WYpRky2L9+bcXG3+u7Oe8gIg5gYiiPQ+9zKCSfWLb74c17Ju3copJ2ckrmfhhS0U
D976Umr9FLpHWaWTxuoyIw+XyWUPc5+fWuC/hnrt2ag9XIbXKuZoHlpnbeUrJA94T/g7NYk468YlohxZU69X614vT4eZsCDwypIzO30K0RTk9mfls/oUdC9zSfqr8OQk
68d7eRIOA7Y5tfGr9TUDy54YA0jDN1abE+Ex3sfHKIRQimQqtE6Xd0vSV5CIutKUY9ltGAZnNc64wjY5t4JegHqs1FrQi/C9hP5IRM4LoISWryZc37BAGn4A1Te6mCAV
giIbrZAfSBfzDYR6nLIJi1BfqacX1prfYN9GRvnq+QmMb1ITSlUaeb2RZfVG78XQYnqLHL+SAegn1g4Gvc2jo16Mzh1Qh1QU+7b7QA0VkEFGG9lWukhbKML9XuGiklfA
et8qeGi62/ZuCN6ooeodZ1goofVIbBdwg/2VAfkk2qs81Sp0+cz0rAO2i/6uthHohjgDcLda82OQVVOTtI9FkSzfRKBtJuREX7h8+eiqgmegIa7Lp33Swf3cLMLA4uhu
0oRizvhnEco9IqWtKECscIgl8w9sXTzzV33y4OO+ugF1y3TBBX1JETQc7Ha1Ngoqkj9UzNxNxOpYtJWp7QZuTMOv+OYDyCIU8WATGeUDWcXsdrS1rnrfhIQztrDITjpO
o+MEsFjcqRro2FMHAiikFPrY2YDejjfW/X0SzJy6fjbvkY+M25nZcu2c+f+k+K43m8EQASkW4oQa7G7rUjBeCKoRvu2tD5kJRdNA5joXxFjW3IbhaVhgUky8xW8vRs14
BIu86hHmQdfRF/lOmDlMyzzlQdeQ+owzABLb0C5WqXNCRnMR7tUMJYWCzk49N/wztqDBgM51VhJvXYSnwn3IYMwbrXjhNJxtWJma13ZDAeWVZnRCx7hfa+PqNPtJl/oo
l9osCSZRrDnFK+eJ337u6MAc94p47mqJerlnVfe/Oy1Q0D6GAqCUc2QOvVChfevvI0k7pScEtTkWTU9+3Ns4KXYxv4E39NNiJCGjIt1Yk7a/3vpjeeZipG4XNf4UcPjz
oW4YR7NseOLCGFsBCQFuU/KgogHIrXQmogvHtJfummyjgFjIbwgy8X9+OQGcaRkvuwaZUAmdIZkS2KqupHZE3L/lf90RiKmaZQkl3x4PUYvBXCSlYANDDqeRpnEt8Hjs
GDxyFBGq/ezegHeKe5QzWw9ZCJtZLWNHWjWNALFutAS+Z/BMkdu4xPxcMWa7CPjWoSWR/gyeWBbfu8+UXaTNdHW/6iaRuZrYWGF9FYl05KNieoscv5IB6CfWDga9zaOj
CjH9J5dB9Llmd77Orbc69MmSLCIsVHIPRjLEIzP9nSQ1nU2W/JfW54NM2rqvVMttsyyrrJ+Qx9di/gw7LO+gaPo5bQjkqgJUWsKB7wgc6GIHmvtRf/Hb2PQX3sgmCAq8
kOiVwGn16Dw5788iaPLGCAhhriFkR4u4vVqS1nAPoD2ayWn/1EJx2Em2c938CLfdR+lRJaNhcNPQFcZfw4Ooh8ePawtMhJ9oR6NJJagIjGYj4ZTvch97T6bUpzS5hhD5
mslp/9RCcdhJtnPd/Ai33UfpUSWjYXDT0BXGX8ODqIcMvZ24aoYIkGAW9rDM0VEx8KsVetiNK2Dfw7HeV1eFz5rJaf/UQnHYSbZz3fwIt92m4fuK4/n36i6QxW0ZDxnH
ReKFB9dgsVlzOduYoY6QY4FZkG+A8zkHXYx7plAANdM6iRe96NdOPtRdLiFScM+kMGVprYnjBymceM4kHmIcfD+QFoSWyE8ODTn5JONswiZEgRvFdNdutYYhyYnb6rds
UdEqD1uvucuPmx4hRVw/5+77tMCwG147cpOzgj9eUoImnXDHcLVp3MtNFlZRh9tImslp/9RCcdhJtnPd/Ai33eVAehQMzkCAgrj8P3CYeirV8tjk9GrlYYzILyXm7KKX
rhR4mjxPGp+WzmA6wEVUDZrJaf/UQnHYSbZz3fwIt90NiQf82HOmcWtiZo93CkH06bgEe2T7FjlK2MgkqKRLfdxpMhCrWoeHN2UN9GZsI6mARZpIgXP4jnYdvreyhXmX
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereGSS1kZpY1PC/5NLBnStY4Pl35V2cz+JKVCCL9yu9bzx5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5XlG9wQXfrGmGmV3iWnGutu81jhkdWPq5sgiw9YEZSGTL7tyVcvkfmA+TQXjH0FLPu0BuIra1yIwu3MMDNistM
tP8SNJzfbqHCElzUSE5Nbg1lea1eGWT0ab1/thS4nP3rFopo4UC9LSNTvoLHMvqXsnSWxMuPZQS7TgMF9GxMaLWQcGyoiXqNTr7WqJYRKZ+LzYKpBdO0R/x68q/7qspl
qYmFzYNpMmhiqdmCEXNyAWc6rqaRkKDMSSkYfWlSqdZ/aGZ91kQHcGcEKUND4qBCJyxMuvdSoPIt83fVz2ok5N05cBunmyR5KMAAondKExEKel0xyJV9ls3Stpb0fCyz
yaGTohwD6C0pLAcihlkcq8YftOCTwQvY8M64dh9zY2A=
`pragma protect end_protected

endmodule
