// ============================================================
// File Name: rx_dpram_768x32_emif.v
// IP core  : ethernet_mac_v2 
// Function : RX memory management
// ============================================================

module cme_ip_rx_dpram_768x32_emif_v3(
        clkw,
        cew,
        aw,
        dw,

        clkr,
        cer,
        ar,
        qr
        );
//protect_encode_begin
`pragma protect begin_protected
`pragma protect version=1
`pragma protect data_block
joqvu!!!dmls<joqvu!!!dfs<joqvu!!!\22;1^!bs<pvuqvu!!\8;1^!rs<!!!!joqvu!!!dmlx<joqvu!!!dfx<joqvu!!!\:;1^!!!bx<joqvu!!!\42;1^!!ex<xjsf!\42;1^!rs`1<xjsf!\42;1^!rs`2<xjsf!\42;1^!rs`3<xjsf!!!!!!!!dfx`1<xjsf!!!!!!!!dfx`2<xjsf!!!!!!!!dfx`3<bttjho!rs!>!)|bs\22;21^-bs\2;1^~!>>!5(i1*!@!rs`1\8;1^!;!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i2*!@!rs`1\26;9^!;!!!!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i3*!@!rs`1\34;27^!;!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i4*!@!rs`1\42;35^!;!!!!!!!!!!!!!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i5*!@!rs`2\8;1^!;!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i6*!@!rs`2\26;9^!;!!!!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i7*!@!rs`2\34;27^!;!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i8*!@!rs`2\42;35^!;!!!!!!!!!!!!!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i9*!@!rs`3\8;1^!;!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(i:*!@!rs`3\26;9^!;!!!!!!!!!!!!!!!)|bs\22;21^-bs\2;1^~!>>!5(ib*!@!rs`3\34;27^!;!!!!!!!!!!!!rs`3\42;35^<!dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s1`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`1*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`1\42;27^*!!!!*<bttjho!dfx`1!>!dfx!'!)bx\:;9^!>>!3(c1*<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s1`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`1*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`1\26;1^*!!!!*<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s2`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`2*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`2\42;27^*!!!!*<
!bttjho!dfx`2!>!dfx!'!)bx\:;9^!>>!3(c2*<
!dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s2`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`2*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`2\26;1^*!!!!*<dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s3`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`3*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`3\42;27^*!!!!*<
!bttjho!dfx`3!>!dfx!'!)bx\:;9^!>>!3(c21*<
!dnf`jq`fnc6l`fui`n6`w4!fnc`jotu`s3`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`3*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\:;3^*-
!/dfs)2(c2*-
!/rs)rs`3\26;1^*!!!!*<
`pragma protect end_protected
//protect_encode_end
endmodule


