//================================================================================
// Copyright (c) 2013 Capital-micro, Inc.(Beijing)  All rights reserved.
//
// Capital-micro, Inc.(Beijing) Confidential.
//
// No part of this code may be reproduced, distributed, transmitted,
// transcribed, stored in a retrieval system, or translated into any
// human or computer language, in any form or by any means, electronic,
// mechanical, magnetic, manual, or otherwise, without the express
// written permission of Capital-micro, Inc.
//
//================================================================================
// Module Description: 
// This is address mapping module for Ethernet MAC IP control interface
// 1. Address mapping for MAC control interface(MCI)
// 2. Address mapping for MAC transmit/receive memory access (Optional)
// 3. Address mapping for MAC transmit/receive memory control (Optional)
//================================================================================
// Revision History :
//     V1.0   2013-03-18  FPGA IP Grp, first created
//     V2.0   2014-04-25  FPGA IP Grp, support EMIF/AHB bus, modify TX/RX
//     memory management   
//     V3.0   2014-12-18  FPGA IP Grp, add eth_mac_core_f_1k.v to support
//     1000M mode
//================================================================================

module hme_ip_ahb2mci_ahb_v3 (
   clk_app_i,
   rst_clk_app_n,
	
   fp0_s_ahb_sel,
   fp0_s_ahb_addr,
   fp0_s_ahb_write,
   fp0_s_ahb_trans,
   fp0_s_ahb_wdata,
   fp0_s_ahb_readyout,
   fp0_s_ahb_rdata,

   irq,            //interrupt
   // MAC Control Interface(MCI)
   mci_val_o,
   mci_addr_o,
   mci_rdwrn_o,
   mci_wdata_o,
   mci_be_o,
   mci_ack_i,
   mci_rdata_i,
   mci_intr_i,
   
   //interface with tr_mem_ctrl      
   rx_len,
   rx_stat,

   clr_rx_mem_empty_stat,
   rx_mem_rd_data,
   rx_mem_rd_ack,
   tx_stat,
   tx_stat_val_i,
   

   tx_mem_0_clr,
   tx_mem_1_clr,

   mci_ctrl,
   tx_mem_wr,
   tx_mem_wr_addr,
   tx_mem_wr_data,
   
   rcv_new_frame_en_rx,
   rcv_new_frame_en_clr_app,
   rx_mem_rd,
   rx_mem_rd_addr,
   frame_rd_over_en_pedge
);

`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
C6aFK2zKQeXwDCX2qf2ZjU/7YrGHyvMzm9DNW1Nh0x+Y+FSps+S5Z0bQy6HvABMh5epxuDJVaxc6OUEcl+WH008rVqeslRKB7/lvkQjRreS6uVPLKzUaHnvlG1EfSP5af/Azg4tOUYcDhh3xVQuPYr608u4a97Xp7nZ8y2K9gNw=
`pragma protect data_block
6so86mxGW2+3cYvx+h5Cenn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3tbSV+HqinCZAllRipm1vxTqyjzqbEZbb7dxi/H6HkJ6
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereLjeLl6YOhMqrFytLZsEyFnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3t45KuzGqziWZsstvq8Dt/MFPHjxKIexqjrqGbhWkIozt3fdWPUxSJL7/HsGftmysnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3szueqiF/XUP+L1nYRC14uH0D9xfughz4sYj0zFHoAFreJwO58fKUl6PMSID/Z6FwuWnPRVETHx+0JWb1oMSh8SE8VFsPafQ03aBKJrO3erQ
AQtt7IdTwpz1H6sEobD+23n964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3hHzJGDIXbd0L+VlwBYBJ8TJVzYt64qzjFnObD4oPxGd
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereR4ERhGbCdav6QRtC0AmqvghpvyhDcTWJgfs4Z0IdDsx5/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t6KVA/McvQg3eOhjeN8DSW77jGaKmgGU3CdTwmeXCU3G+EQat6CuWI1sd4T/rMMxelrBihypB8MW+yCGVa3tDA0
jfKFQQgUt1Un511RVJvnYe0TrdznDtCXjr1MVar9OM1mVHEVWrjRI8NnPi8bPzHLr7+Xbbe2wKCPDv7hh2ianedoPA7MDZG3UmcjY/lD2F55/euKxkcULP0LTdZTgere
9W9wqYaeNf/IMTNJU2zWK5rJaf/UQnHYSbZz3fwIt92kGX5PRo96zeogAmEU4V2VQboXcX5iSPmoQ318BSNdhn7DdPj44TkCrW9Kulahfc3kKyqlihsEDSR+CqCXSHot
awYocqQfDFvsghlWt7QwNHIoFv+yh64xHZHuNLNbs06ayWn/1EJx2Em2c938CLfdYSB+dWPYrmhFtGY4Y7Gd8ntf7BcdYXqeScS3UKj2/I15/euKxkcULP0LTdZTgere
LGFWj/NsiJOnSuaOOwUMVemCnBcT0x+t9Nl+hQwsxyTwQr32Cu7B/iQjVTfoozxcgj4thrLMZzhuSV3zTZItGufJgFROjgf72XaxM7eSdx15/euKxkcULP0LTdZTgere
hIAuAV2Yc0v1Kq83azc8/z5+/uStayjc0uWse0YEnwZ5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t7xnlyCEMyolv9C+sUwOTaL
cFW7o0jCCghShJkpxkyfrHn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3hpp/L2zeaLgckMxIONqyhWPxDA/cpxj4qpQGYvt10Tc
ef3risZHFCz9C03WU4Hq3ub0xgG1vZYUbjO4Ri6BhXOayWn/1EJx2Em2c938CLfdXdx2IEYsYU2Zd8VLQjllTUMw4zOswa52DXbF4DDxJ+tI3QhO3YjbLGG8jp+8YjAH
o+b8XKts76nQWqvbCCYrA43oZMx21C8yshYvm8Tf1MLmy47jWEqj23E+y7mYJex6ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
A1olyXfP6WWXB3efTW/fXQVkx+QwcRA+3X2GtmpI8AeQje4FXjJpjkQtkVQpz6P3OOgvok0mtjgapBTvc5ynm3n964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3mKPPszTlq8JNNyCnPKmQzFRHwarvP+uRzlPY4bk4+BKozba44PbADasIfWERMWAIHdadxFlhcwAaK3UvxNBEMyFsxe9kI6hCLfQDTeWxmRw
XssnmldPLyaLwVLT/Ox9mvzMSzcbMUCZA0EOwlCSqCAzk4hve++dKDnyVp78hUEqWJATxTYkJ5Bh6Ljfy3HJlm1EgUabgkK98BMurn5OPwqoEkzQ4vSPEPBopLfM/9Al
Nf5Wp3gE2Q5F9L8FJ97VSRSvYp2RgD25FascNnOwxGgwyGH0Nyf1No+1tq3R+tVKDx9iNjPLOLDuJ+EYrphIeODRrMEbQDd3cID3tkNnjI4wWCEQ+ND9y9WozszkCWuI
pxeevPef4x0g+0747ML9nmzHJy3eWd1MZ6CMf9mDoYhdSs5546R0i3q/ZHnd3TJ6wwk+KCsa6N6I0CSsxfThKm3vizlao2121Pndvu0cAARYzbhs2gmfvhAPkjGhwOY7
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereV5RvcEF36xphpld4lpxrrcBqdvZbGjxqx/wY5Acvw59MNZTVeicENM3mi0YbYj4v
kj3EI+HYpijsKxL2bgYmMsEjMDe7cB1twShSmyf7QSt5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5U2mOCle7OJm+bad16xzSq
C8tSOY+Bq4AilXkZUHa2NVb+0HaVWpu+oJdhaiKMAcE/Kz6BRWcyEH90OAdS8PKZWQv6+REik4bJjiZKwFEhBqQG17tHMQJnIgObjgEY59SKJUao63TNrEVGGNgR19s9
c6EIUiGR/rYjHLGG9SLkm1+AvvsxaIMLCTktMUXnADNlnZO1fn2TlwW3HKvaTIJ3m1SFyaCmy0ig+/jIQvrfDGV0QgTd86ejiIex1wAtDlQTZcHMSxkStDY3BWA2YAoy
jeiZxI87MksNY7BaNNyjbtBjSXf74KqTnoa6meCygVOoHBwoOOrSxajl2vCFvA4mEm888E4B5OP4z7yPX6A3ONuKh/nhXiLFCKb/PPebpx1UMC3fpUd7GlRkdX05rAHR
98zeP5CqJfa2ivuzciO8gYUlLWdz84vLkwA2dJwVpLWGFT9wA2cahqRkm7cb1t4zMTELeY6hcOrceRa4Os02sOBguB9QXYHZ0wqi/NyCHrHlydZrzILC16EE5VP3ZjD1
2cPhT+fdcoM4LdBlIGF8Onn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3leUb3BBd+saYaZXeJaca63Aanb2Wxo8asf8GOQHL8Of
gP6tLCiCQKBNMy1INF8BPjg95CTPQZCNKADv7qJAjdQjMD/TczAgzeenoUyQCjzref3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
+i74+TopZ39QmB5sihC7e4agXpjGXKJ5imVTGF5Rba6UnSMryW4NK5KZW6rbC2450p0H5WbJPsTAEGXu37AKAYqueKFn7IDiJTLkbPywcxRaVoBiXga29qOtNGELuFi8
q65b3Y/QBfsbWoRgYBSYFC9Pzv5LFBbMRB0cKNiZmqQOtQR6Zl13TCn9O+D9LyVK+sFhmQaDVw2MPiAv0PDSCIHTmJP/xEvXRLUXcJUiTk5u7MRtUY/p1cVJDiVJnG3F
O5oFXDuswKi+eC1Gtn4PhHn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3ma/Vk6+5DbReoUEDAISTOWXMD3otA7vTd4NGZROpPZd
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereV5RvcEF36xphpld4lpxrrRBtJ9TbdMwYV++1UDC7rq7+YOVWAj5DmT3QDABCwO1L
bZIIpp1OVoC/N2+b3Oz61Hn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3gCDoYn1Gnh0W14LaEj7zB0hlJvXCu9dW20YXJ24Rj0k
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereV9QT+hnGPjc9GUi7n00Ode60n4wYcPkUtvifA5QLXNwR3HPilNhIBymOLMfleHuF
2TdT3Y3Yjrq6HNHktrEMWYV2G5Z8VUIx2C8ImEXrlmubuSntM9K6SZYERNKbXxAQj+fzP5MIIXAP/GKb+P8HLkWmo4YFycKQmEdt1z0WhtWtpRtAgsxtJ7SSx2YVJBJ/
yK3/ftXIbgsKmWc9HSaK/iGxlwSuYIzGPIzpV7b629i5iFdp3HIuMHtbdr6wVVrplDSlWnx1RGgzzAxJzU0MaZ6xaxU12L3evtm4sF7hjNOHE0aI1OJ3/WKpB51PGJbz
3+Bn6QJuqN3ZZ6KwZ+UdCXn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3vJ+wniVMsZPbzYfue8TAqZ5srpOJMvGu9tx+vwp8HcF
81ZCbbLcXPITHG4UybLxUCF0c3Szs7VbhYaMLFdCGPt5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5J79SH3+X8M1tH1wQfoNko
jsTV9y2GvFXIZmA6pF0VrWY1SL0QGszrtFaNzNTzj+1ev3bVYpOe7nWwo/x7C5M51w8wl0U8vpw40JfspsV8HwDZqywZarIzKT91IwO/7pId36LYEZHQxiSbwWS9y931
O9W+qMj/j0BieTEfARrbLyR2UbmbwJjhTu8qVXF/83Z9+7qzydS+ymhDVkUll+CFlf/2AXL/rENn1udcpoV5HxiKAlFj8CEisSj/TGng/QGDIqojtL7EMAa+Sf9WesJM
OJKx674bMVjaKnMK14QHhMmE6Iu+aVlQqTml02NO1+XxzNcECGL+7+Zh0MfObFpoNrYYWtKbGuZxGUxjNAtVC+jiWpe37mCsd+Vt9j9E4/xNUEkT9jq1d9BFYJGbiuC9
VlyhqPCg0QSfBF/8W3NmpoMuDym6eI40tXIfpBsTddQXuR3+P45255UB2/xrWDYjJrMLHpHxNJuy4b795XPQ8s1iT/FCVAMBJhHeOFOkA6eIRqsVTTrdR02/BArqsU98
XQvDSiCn1sYgZoMXB2UgcfF8KPrzG4Nr6O1WmiztWmsRxC3OLpaDoksgBXhnx5Zp+3SUPvI9le3bCFO3ZMXWOeNouu1aFNsBMhYWgLCwe917tT4OJz1e955Wv77jO1FO
QEBovxq19XGL2iMtfe07jcE+OBvMkg6h5KsXGMvY4RhSQZ5v8BEMdbolQ8IA3txDwLghZgPDslTf4W58nwBOKx95tl2wChGLWs/Akzr5MZVnkA+AmNaVJ2xhGDnQaKKe
ia3oupnQgA2OmwZYp6qLhHn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3k023oXTPcOko7Gt/929+t/tThAtJf6BCXeIx8MDPZMP
HBQBo79XkqTXkfLh3jgmmhMb7V6FILzkKA5jgQKCNPXFAAyXAfZ1INfF31EbUmv3ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
JTohbGPorE2HXOHo+u5JlGY4VwiH1fK/vakyCqtom6NvyzBX59/9AptjscX2cUY3vmIpl1r7NPycD93o/oQWUbRGhk4HnQR+6Oqc9zteSW8tykA/6eABffq5WGp0RdYK
PJsIo6GfcfbnHyAmJI471KkkQ+gQdCvAqIzfqFaGiz+SrfCnRx0mfzJkVwzRxHOtvVCkm40MXMcv0AU34oqaogWkgWg7/PpIL2ufxHd7DWcAdclvVOQyIBxcRTFnb2lz
65rIdDBihOLANS1oPQpBs2vR3RgoHwVOuA6OgWIEdOxVHi6Ujw5doG7h9tFsBjXmT/FZB+oa7o3yJqA1YHZMwazzyyz9RW8QkcYCH+J2YhQRXe7f2sSETWERWv+ZAiCj
CDo3Op8Grcif6YKNc2lZyDWy4bfAMGr7LACmoYsDkaKfzH2jjgsEVRnaiQB6JaM11M2XM1BdV5sMvx9eNgH/a7PEpSO2lyF1D3Cyco1ZnL/+UcefQ24/56gTSlY8Gc7n
e23g0mIkYiWqkD+/J0xQZKi///+sd7BoEJM+a7mzJCsS0q8/MWLVBZoRHXlj8Jk+BW5xeX/chsk4X32rTgXJ7aKbx8qruMNgxUZEjtOQgU5wHh21oYZ1GZJklN+TNOjs
L1esuf/usl2uf5N2vHqmAyQtUXyrb6kX6LKLtPaGNqCNfzYvb0p/Ioco3zqzWjdCg9SSdRRm2pK5QBJD9bjYQgQRlVCAcyVsw5Rupb8YeWuuZSVPPLt/m1IHsrON6O7o
5VSJhALWSzR6e9MiZ6fbfHn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3kqSpcDiJGQxVazosTEidf4Q1kI+4gUFc+XCIiVMsHiR
J+Ur/ezRrxoRrRe7gMA4gXn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3jqbM21w4nooYPHghirkBEJCeHP689Ex7rmPB6sExH3u
gTZx7bTfLJvohMoqH2ZP23w2wx8M/qefJESwEoSnSxlblfARpTvOx4W5138sClhriZaIJM6lCmNImt0wrVGhfVpyXt0HT9vRGlpU8KOOQmjBASRSXZuL0wiTOSGRr2EH
467TzyQpIWVLy7VLzH8j0iDbFRQLGxsoRRidAWAfLllSfIAS5TWJKSI3WTFyq93EnpGpW8HhTmLjC5UpmC1Nbdu1/GmvZRKwAi9b+iEq00T9UsSyKxcvb7lzbrQtQ5Wu
Zf2GICOSvsTt/WvnDQxZktFLFHCV4BpzRZ9IyWM/jF4zVCPI/GIDnQJprwvPz3uASqiOvl4loAC8630wZBP3iXwnWzyLQOKdyYIFw7fAUL637Tf9LesEUoIt58Bd//O6
uOzuJTr2xCg2H3bJPiM+wnjizfhH/6SnHyZKcNg/yPLlgZVSm0TQiNUsHhSf/1T1ib26SFXCNFCbQMIaVrR8aqSEDvVsRuzBbxaAVOu711v9sjAgPbPU53WFSfrArLTs
fADWXBMuG3hf8u6IEuREX2go7eCXN15YIig9AX4sk9TIT96XiCJufEfrOBEobeFVhNL4QmsYA9SCc9jYqPMQNShCdzODtAM9mKf4SJRSEGVW7nfsYqmXp3Y6yueGUSgC
io8wypo3GQGkd3qh8FJZ+rCL+bztWQ391wrkwmkIdhp/ezE5GFaJE0pEkC+bXztvaHkb65Anv4UUEqYJctp4P4r20uOR72IzFsdjgXyCSGjgxEheqgzq3aQ+qbJvnPoK
8BndxWmXbhROhzV5dJcSR8CwNF/YKr9VaAMtsWC5mn7i1ecrLJEKAlZjChwLIR6XZhUIuVFla9O7/XLyR5fdeNt/OEpYE1KcsR1cVbkBj7Oz9NBFkS6aNRvfWNzOB1Bp
hcUWE6a5gXutgcmHRpl08Im3rNpMNUBNZs2UglaVJBVB2oIIIGDl2Rsuyl4DIOo5v3LpShHOQL/znZuSzrHTXbSokJJfR3bmdswLCb11hKKC12BZczv/nh2Q+Ij945+C
dn658w4qzP3w+yqGcLkgjevhn9nLVV0NVjZHoRuabjfi5HwNMFDOzijeV1/U2HpozNPu79Hdz/FRxTBUJVv2TwL4F7pRdO5cKo8OxIsfO40yjYAHBeNIqZuHhgtmtvn5
/ZFMF9WQ9hcbGmVDR4dc5HF7goebsYBqtNNqTLe/d3P+c2gRRQmunSv1KOEhebizoexcGP2wRfNPo8b010BcMhIH+849PG+tgqezSeyQToEK7gmfyGXjdFF4YiKJ5K3R
DeSaIAvfcWs1h1ZwXxU2EEoUr4iWYzc76s44bTZxYw/gGgUJqePN9NuBXCJHdpVOcEcYZKcVPBk2QKnL51OjhCUUYqolgcz03AnqfHXS+DpQqn74FyEplTvsQY9TZgdn
DQrLQI6aWX3AwoUku+nId3HdiPqmYzxlA90urkIcK5Ctnc9TwjPG1PwHE3iQjcIW7zZj8mMFuV+9n3ygHrPAbNntQXa15FgZfoeJs2ikqfSUNTyY3SZwFLvcN6m3+40x
cTBab+mMAheQtfdjK1pg2sLq+KVlT4qOPQ3SdavxIEd5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t7OwMjt93CCpRgU7eE8EWi4
pWXjXU6Vfeh0eyiWKBQsMHn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3leUb3BBd+saYaZXeJaca63Jny/DY0uI9r4hag9RYX98
OqceS1yEwLIm45uGYQlIpS5aRIka8SbvcwwaCs35eeJ9R2qPSQEvAT4yP+2a1XZ39Bei2J23jKNDylSrks+RLDsw+PGzgnY348/WzVgbZHqRzTIeeuTPxJn5QwTlCchu
PVWdn8Xq9Z+EiWuO4otG1CIEeBehQYkqzlfL4MJ5wHdCUiKaeOLsUR5TWY07bc59PCl5Va9LPPDH6fTVcxQEkNDfSaWvQ4B+2SHxI6DSI0GaNldEzjciJbd0KRE5DtjP
q0eGhC9OaZg1tHbNg+wZrqpYVSSVB8VTvFN0/c7WjfoudR35C5SNkS+ESiFAxdJpLggltc1R6dRpzMgst/dLGGBu1OPioxNp1BVU24eUp0YTpX1VYyl3hXU1kPhhOrL0
a4Tx6vqzc9uEOR5UgXpCuAbeSf6o2YV5JWjcplH1WhyE0vhCaxgD1IJz2Nio8xA15EUWFiGO8G9tUu1/9mEOkEJeiIAmXYIhFSxQ5IK1ywQIrfGnfXf3bxfUjVWmzDUB
jS/w83if/8N5xOMizwaFVx10tgRcnGNagLN65QmNO6WVeTm2x2W9j1IJYuhzyCx9abBQVpmYaa2rerosJ74YdyHZgC933AzigTzGcqdbXXBxsDRq6bNdVVza63jENPAg
IW40k9xu2HCkNyv1IHgYsAkVnxBiNQ4uDsLcPuueXewJ/qlLamFsqIwX7sWTTckt4nS+uhczsgwY7HMyLoLPa65cZ36xSo0K5TYjqZEG6Acd6Joo3F/jJmWJEhXNVdt8
mRs9yRC3Kb0hNOeopEpKXPf1SDjQ0avq8PsjPDlrq8GlHFH5+h+i3TL28ybyKjRTQqF2fLytTQBRqQO6DDmA/p3e8IZ0w8XP7N4qnUrC1MlFGHvXvZA+KUHFY5JXbd6h
1ll2i368HqRWrR5tqv/27CzfRKBtJuREX7h8+eiqgmegIa7Lp33Swf3cLMLA4uhu0oRizvhnEco9IqWtKECscHHbRL0aJXjDaj/rEMFg+/B+MfSIv6lyhYVA6DmL3AGx
Oy6/Rq92PzlABLYouRXbbqPGJwlAGzJmle4df4MBPHH49277CZsTyGcosC//WWLfnarotSvxhWHsxpp2g0a1cDEe/5ux7IJ60mmHhTZOqFft8727uV7QM+WPTa80FPXQ
FNmeQz30rkSADml2bqp7jOJN14nFid4FG5XkvmYuvVgNrEKbE+PV3jnumpq/lmEb7/vatlzq1CKX4FNamHFwroFNLeEiTq6mLNOg5eDXl4tq5LtiwFzRpIWDt+iAHjKM
kVK0eqZ1yE8xFoN7nzTwieAbI7wBvWlolh8R8rzIRl9P4c34T7UjuQjn83y9lX+imLES2qcZ1KgVOi/vZgi66+bHRLyD8vC4lSnQHWoC30NNOMCQD4D7bydr4NcrsVfj
olk9dyBMQ+adiVEJhV+iJVR8Tr60eMTizIWFTzRJnXzZT18+7D2q0hIK545bH67pXBjoDRCebEw0K0h3qmfAhoY4A3C3WvNjkFVTk7SPRZEs30SgbSbkRF+4fPnoqoJn
oCGuy6d90sH93CzCwOLobtKEYs74ZxHKPSKlrShArHBenc2VUxKrz6oEkqsCjoEEX32hJopJ2qTwSa5wk1ZC4227AAel4SwYgCliXbpn+hu4gpq1o8LZ6EbV4w4XOEYh
7fOLdNcn6B3uyLKEHx54Tnw2wx8M/qefJESwEoSnSxnyoKW3texQEnOlOVDtCPaogJrFf4m74AWImR0hCA4U2QeJr2vIQ9FOCXj4kTlwzNNbqbLGehBkkOX7lpx/sCoB
p9snHgtHT1nWx4wf93r2kylckX0Ct7GQ/mgE3dxmTUn+9/qVQPzxfOxeDrGwjY/dnIa9yKvRKRIW07lRB2BunZWkw+mQByZzMgFjdxxOcxoQu66ehtl2fqWm9RmUKrrS
dKWXWBSIm8zc/fcwTl0esJ6xxJTMyby4SuY/IyIRi0cHIPf5Heo5FvsmJBIVUI0rPNWSL8utZMrqWw1w60iwLf2igJqMbsc42ifkdFVObbpkxfJIOs6elmg8nP1A3gjD
yy1XnJvEcmRYxgQDT3o9HFDPOHyNeTBYipdHEI9a3Ku2L8NROgbDPmK6G7Cjn9Hm4+VvGe6rtYg1HmQQA1DsAvH6h8mHKSz1B5JMeYtkbpXkKNJuV3sss44CN4rMmf80
WYpRky2L9+bcXG3+u7Oe8kUmh36c4MlOkCV2iUQTUbLumtITw+MenFmUhFDwEtglfW1v+c/1zgiRf72wIYsvxXJWi/7spqZLkdKUx1t1VMbn5JjPfW1pBUaSQRfq4+sS
syAJgBa/BRB1nMWV/2zB57SHQzIcmdos+725d1gF17Whh1oFthKSiPIVSoxZ6cb9mVmhr/M/i2HBvHvfUJuGY20TgCWfJ/wAnEDaC7buh4aWMg8I/R9ubMrigUXcsOdy
WpZfs3M7SFj1/UfOb9pSuV/3b4SCJ+R6hHPSBztOWnEyT9XHTRfO9hBTsMJ8/b8Ec9IKcOr5GZyUNbf9DzJznWCerPo7q9SipeaPyBKB7Riyl3urMnCEwl9sUsgS0YiL
wA1sB9NV708BjQEKnMde1c0YAe5ERNB5XZE0RKncWaQA4/bpGF0sS/KaSfIlEm2NiuwozHJCASzK7M5TpJeLhuUffqz8eO3RSArMST8/vwnU+3i+C+ZNbZs33NeiU/Pl
HdAHkJ8ohXu9xMc9VQJRkbH2+Y7NSn9ZRMMCL/m8+rpAk04NNuwPkGrYUvw3uk/UdOO6wWSObWwFxpaPtaU7RapdiYbCTMLeD5GkK06/fFpGat8zcz8PtJ3gBx7chdUC
sphtLhdFJzwOhMd6TzXqKJEMNHjwK/TfCrIgimTQpd035NODenyZYg05Ap7GYrLVthwXHV9bWcOspvCYxL5asaYksUZAhnRSLnYIfzYAuwDhZZmbwA7voRyD3BMcapby
OsBIbOXQVLRAv/IiZpmynQVZFRK4ZoT8a6FcmNYyNBwjd4YEUbxRLiaNqN/ckbzP257xtiDREYqzbyhlVwgMHdwRAu6Bf1zLCnEQJH/lTZpQB3EoTOnYtQmErQvUoq8E
C2YmkNSryxCPJ8/3JCVQcI/mFBUpfRPlEYhaABPk0brXt4gV4W54Uclm+tZt5yKxtkrng5ZwZXNaFk8N1hY7YJY0VGGoaJzElea9BBpNuFrMjRYnxbARNNtk+iVwmHAI
6hGckDRwYKtZdxdTPTGG13U49F8/hVJGfqR+/x15tismR5WWbOzXnzunngXkq5r07M58OvuGitQizSh22rzi6yY6pIvTmjfe4hsxcm2Qu6my+aR6H/+m43B9iZv1ywiD
3tNRdtE3k2/Q529OmflCPHDWy/lnmacEfREPJE9CD/A4COM6xoAXG4zSOs4qks/XBUGZMOLkiwBnxeLbJe7nMsOiwdCnnQqTo9x9IO9MP7wQES5cy3ybmVhEakap/eNF
L3TVDqt8XKfiAnV4apvfDw3b3zkDLIjmOkZIIf4MPqmO1AGsWvh+pPgafPkLZd+6ETeV7X6ZrmZeK5kKJOY75vFqH6CuRdoDbVtzJuKynuhgm8mifPGWo5DMp81YiyLr
VIB6ORZMgdxu7frB6GWB3lLI1x8+x4Gc3M5uEzrXeAGRVw+q2G7u/cnFDltVb6k7sxZ01yTdd5hbmTr/ie47LjLVfEpYtw847B/AryvBmbGyasAGHJiyLfyGmWtb2Vbt
0BdEPzzDQk4R0aeWQ47SC08vcB3CxI1DEbRnq24EQRpUKt2BUGUeIT1t/DM1GSrKlWOsVoKcTjUAAm9l/hvIJWIcriS5ddDwUNb7kFm78UgS5snzjkNTfwv8vnK/Cq8b
fW1v+c/1zgiRf72wIYsvxbSF0syRcZkX6RVux+8e7giNAzkhKqOzJIUpJ6KaKAnwTXmHr5auratDpE8AQ4VBUw+tfWlMMV9fNB9knho+KZ1EPF/KArXPU/8U4vsV+J0s
5gRnkq2wlHjnIaeDlqLnEOXojXvmdM7rDTnFcpCItAMr0nDzU9qNd+OXkC8m+f68L3VRiA2P4RfqO7zmBzn+3YZsOVA8issbREBxjwYZLEfiiZdVsAaNefwgoScTQ02R
e3kt/qPj/iS0TfSLlDPjB0oIr3IAkv6Hh34K1dId6UaayWn/1EJx2Em2c938CLfdTrdbsbjUc/NbeSlwJMqDVNWjQ2TcBfpF/mLVkFMmWt+aDo4lBB54CWPzgTWhInlj
4EAqJTfmLivpGZ9Q9JFkYJrJaf/UQnHYSbZz3fwIt91FDOmevch0lGe9hPpwI6B95BU/38O9tVDAR1+pdUU7zZvMtqb+W50kdq+0CBqLJX3ddJasYAugAQhuq9KtzfwU
mslp/9RCcdhJtnPd/Ai33ecK+URBqtbpzYPx5OeEeBmwQteCZ9U8ed7tNxkVN1tsYutXsBejWIenw6XSYch7py/KaU+zFFYd1ofx43VCsr8tW0mzTjKLbNdBcQ/0eEk+
hex3QnELA/P6u0QOBQ5fjnu7lHx99sw6kFcWWzc+Xwo8tWc4kUCBF5DPtGhLYsBvLNH69pJjAIW/KiE7dteP92CHEH2PVjc+uj+l7UPrIZRN183v4+/FpjY2AVvsagCN
wM4ESfwbVU1XoLqMFaNLrtxdnOOVkeCX6uA/Dh2o328ohEQDAtWTD/ujLRjbNUZcomUqodQTqf0dV0AptDwybiaNOAC9+ScnZkjRtS4uiF28vDJTgAwEguPMYvcnvcNQ
SglyKuqa2dJ05AVMUOYdL7MoBUq6Lg/njyrSlAqJ5deayWn/1EJx2Em2c938CLfd27CdSxwXM2d5URARvZj/V3n964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3mpHuPJPMj7FzmMEKoda+L9AWQirmr7R5DjNlYowLgXpP41SmRErNq3A1ImMusmnCnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3vYs8QshIAq2193OrBpC1MZ/gw3Kjb8W2BahmBvmhFLPF7W/9+gj7127ZEm6rLF1VnWaR85TNHjt5rJ9Izds8PKyppEkVOmDfBx57c/cpF3R
iWGkdEpVOHnpKtRxDXcBw+d1y72DV7SHk8WftLH6cGplQR+iPwGewckQb3Dira06ohPGfFy6elIaQV1xPsKl8NPmb0zckxkQA5SGk5aJMVPtta/M/aPv5rWjus2JS9s4
5ffYsCgZSJ1tq+foqtZV32XyBW5xYbX9dttLL2UdG7XYdoVCGXmzWCN3UcxOK+rcLDRJdY2R/zewbhWDajGtJI+acKgThl5Qr0kbJATjhQgBMp3l5ypEqSgDrAr3tDVU
qpn4g0Mtrw32r4QslRMDfMsJOpqDvXx9wb0zuo6MJqmUFJgufJRz3apMmWoC/11Utq0Tu2vkjLOLRMmjPbRA25ba9tkNTX3Itc4JgToQ9/nr9YFSyOmWd9Lx7626u8a9
0uPZSN6SGgJYSADpiHY8EGMiETtgeaN/CtwYea5GcTPyqOpvdlKkQ6U16E7n+GApu8P1RJOlNam8IxJZcjTRpRaVRfKmrum8IMVOIt/NY3+4mzEhoJcKutucXmQO1lK8
g2aTq9Aks2PlfL/Iob22yyjGIAgo7/g/8lF8gwg4/hxmAvw135Ejk31u4IlYfmllcrmWtug+u4OsMkQHP/ZI3At7NtI1SzJHnN8qZfU8RuuwDEKtwBP80tlhPN4kI9su
HRDC1K/UqjtDVay2GpzlhS4Mxcbjdxc2sdWtsF5LQk8lWJvLiTSRjPW7xfQQo4/Ukc5ZnoPjwKAbTw6brY5nDk058R6fzqlieNzh44bBUumsx+hXtKTDP/8ra12Pzw/o
2DcOvigL3sbb7H4m+8jF3Z9KFL1LESFjR3TlYRryF/ynJ6Q2nTBgalC9HFOFFf8t0wmydHZv3W4dikwJlyGo+OW7F/MVHSwgCjAilZuotK9x3Yj6pmM8ZQPdLq5CHCuQ
YhDjSeI3pHzwqqQZxsaYjhzfB+ftXdG9/wKG3myM6D46ZcEOcvWVLo2e5s6bG+uTrjeNZZy3W9SqtAGGTUJH1YEbtlADBcBjq0fe2MMNXBObT9Xd4Nr5nZ1Qsl1Agv/r
ef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgereZxi1aHSonvBg8Gzr6L4pKsMgwXBxxG/NzmfoYt9SDmkNmOeS24aV7Nw4HFbXU5/d
mfH3Nlvd1EC8S8zNf/qx+GevpSnQ6K7ozlxRBtz7nH95/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t72LPELISAKttfdzqwaQtTG
f4MNyo2/FtgWoZgb5oRSzxe1v/foI+9du2RJuqyxdVZ1mkfOUzR47eayfSM3bPDysqaRJFTpg3wcee3P3KRd0YlhpHRKVTh56SrUcQ13AcPndcu9g1e0h5PFn7Sx+nBq
ZUEfoj8BnsHJEG9w4q2tOtHH64wgVPLLtYnFjcRNUN++XwDusTkhXGVih6tdn8aWYk1r8/rUY37pkL+REr2JLd1vGVruwbwD3kDvMe/K+4Rc0uIKgE/P77HsSzDQY0lz
5kOlv/HnW45Zd5Bmx7pNbfmpsda2zkh+0FjlRek0dnsiW2eWlZgMX04GSH2mmTE3ff6ht/G/E6rouN+qDYGOvxQwf0T8e4yTd0ZN9zBDyTPvim3wpiaXWHfPorg3XhqB
tONUATi+7BEw9og+cNRxdXnIgcL6pdwm1F5Y/xVoypUBRm1R32yf59dm3W8/L8E/7/vatlzq1CKX4FNamHFwroFNLeEiTq6mLNOg5eDXl4tq5LtiwFzRpIWDt+iAHjKM
/8EduTizEPI4Ids2WkI5dBDQrf6o+OJvCILtbjf3IxPJDlSVyFiW3yPGJVUdjkePXtNBcSczIHxHRrezn/eqbsE0KW0UkayCzgUrFVKjl2OClXfiiHV/3Ue3WZNkRXXG
w5n6tBAnKAkVg7MpaIuGnzLBRtb5Ox2zlU25m7pe8XsVVBPjcWJ6R+duvFNcaFgEX9O77A4UD3Xewdhjm7W4X48Z4DCdaEvafhB/C0bt4L4ew+jR5B/DfNwjEDVKFyla
5zcgcXmYty1MeYucH3n0bWavQfnSAoacvqwHpnQPo6hj2W0YBmc1zrjCNjm3gl6AeqzUWtCL8L2E/khEzgughLG8d6zOIJ3JPhy6ggVXwdyyl3urMnCEwl9sUsgS0YiL
MVDzosjRnKtBMExSJdK6lt4/lvKdrLQXO4X9EABpzRFf2Jv+zvtiaIppVof16ohugqNkdh51au7S69HDGEihCSLdsMftvDZ2SCuGde4Ke0F4vD6+UczGm97nT09DzHWh
cEAZnapYZLkHyp/XHYi2xF1SRtrRYON9Lx6UKogsfSc4CqZ9RRfeGwRFo+wu8U+Qo8MO7PDSr6MI5ShAfOmnukVupUom3guUco5dCEkKj1QKlPzNDOKwV4UUSdLzy4IA
/+Kkplm3QPKWi+PrARer9rLmBihySyzfZEYryQFaIcAc3wfn7V3Rvf8Cht5sjOg+MVDzosjRnKtBMExSJdK6lprLUPZ9xwnWfVxZ/oWcAPhl2ZxjT+8dJEk03TAjfjOQ
j/q6pilzKrmIMUD1pp4DWskOVJXIWJbfI8YlVR2OR49WvgOoJXR6yz8RGOlYF45BdYWMGoC+2SoSP4tyJaiTyqGtPpq3CJBWff/Mw3I+MV5OqWw9Htp5VKntKj4+W8Hh
rzSLu02HUlLv0Nto2n5Y49gDfjw7S46gWeBpjbtEbMZ719RFMcaDyls8yNAL9VKIBHKSBIjVecLdS3QSaREwQZ6gf0fMwPkopT00zB2zwtBimMquPVWg46w942Ocb9bE
TLWGP5I4NUgyRkkFInDvdLNpNSIorZId8S/b3FB60O6b3BA4k6gaER9i483f5mINef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ilQPzHL0IN3joY3jfA0lu02zfjpn2VbP24whqlQNIPvA10Aq/h1AD3rZoKzfz2BqhPakg8a7UqCNbmt2cesOCnn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3sv1Clcnm8Ur53wYECStDIrP3bx+O7Se4Xo5wa/Y8wWKbvdlNPm14kak7h2mUBMV5ZXNawJ0KAUsn/9CxbnKdeptmV6WIjxFyCG9LjYDgTKN
Tdl8bbmo1ENvn0W+97PhQDrPYCvAKDCIPh0h99FVqZRC0qasSL3CWk2zzru2AJWeUkzEEJPy9OqdSU4fxXAAjhdncsPR7GR8lRI7KI2wGJnCheJxTEHTYHFeFfkZkBD4
6nyYlQ5u8uew6937FTD/tafbJx4LR09Z1seMH/d69pMpXJF9ArexkP5oBN3cZk1J/vf6lUD88XzsXg6xsI2P3ZyGvcir0SkSFtO5UQdgbp2VpMPpkAcmczIBY3ccTnMa
J+lgO/Qs7UTa+qWEVsdPao9p5a+UFl4TALjX3/DLSAWIxEVeKxJdNppxHvzfk1Zj5JSdr/bnYJkz4BUYGlBmEC91UYgNj+EX6ju85gc5/t0yi16tIPRnlwdWMd6D6AHn
nILPFl5Hj76hDnco+8lUbkcHtMpzIgSty69NitbP4tp57XZJfQ4qt3wLI7dtMrGs/7kybCVI+3zkYtIyOVaY53+DDcqNvxbYFqGYG+aEUs8Xtb/36CPvXbtkSbqssXVW
7+ktrBWVDKEPfTmVtxc90u/72rZc6tQil+BTWphxcK6BTS3hIk6upizToOXg15eLauS7YsBc0aSFg7fogB4yjP/BHbk4sxDyOCHbNlpCOXSBFlkFx/3+0yn8ohLS8omE
JotFarbKp7G07DCSINNH/HxpfeG7I07PiJQexTYb85mG1C2Y6ESsH3CVE6vce/6P2kk5oFbFuul0X03Tj9yhxJ75CvNL1+5wlHotOQqMbtDo8hSmg1oCmiUPae4C8+Kg
viccvvCLUEq3yZ50SXjo0PpwL5Zj6yHSB8IzRFqARGsywUbW+Tsds5VNuZu6XvF7p9snHgtHT1nWx4wf93r2kylckX0Ct7GQ/mgE3dxmTUn+9/qVQPzxfOxeDrGwjY/d
rUp5+TB8OEDzmFUii5RazMk6gX7ForwbmXnyxf2ahpfaLzYc0YZ5VbB8ZA7eY3He4WKOY1BPG8g84x/fL8F/md9tmvv6eBEfUCwTAR+MV4ojxLMr5SfH6164UyD8qfkz
tqmbQmPatbjH+GzWb2gk/VhrBiT1qwStuEneAwAkQgFd6yT/fN8IY28aheYANtbLrpilOpB52Lkf4EBPZHB6ASPF3bjF/WimU0oCCJtX3/SH8yWr8ApWtw57a5NwbA02
iEYHFErUNXSZA+hqWRT0S4Y4A3C3WvNjkFVTk7SPRZEs30SgbSbkRF+4fPnoqoJnoCGuy6d90sH93CzCwOLobqe8yKDh+qWBDonlitJDBF4hezaLC153XcyfPHvNWxbM
hVOto+nH1NMCYY3RGnXToJflkIkZVMNlEHU/esIy79YytMswt2DpdvopckJEncmB3QhVutmOZOU6F/DHUQfrSfn9cMpzPfrbl8iDFRkNY9MaSqL2eRbQgsBlIcqXfWuS
Us2dyLiNDK4lFV5lYGtOz7dwGIUN4UxB2Fz7lKxYduRnMSr6PTKze0alVgMog77CrYsHq5dgtURRYnR+GUnltTarKYGCCd7DPwYsrZ4B0+yxShf7dy3jv6BhiAuuSLOQ
8zqLgQnti/9ACc+cwUerJa2LB6uXYLVEUWJ0fhlJ5bVZ2wjiNjXtQH64ZqKMP+OdeB1l4vwBxjoQr7j/W/Sh5+/72rZc6tQil+BTWphxcK6BTS3hIk6upizToOXg15eL
auS7YsBc0aSFg7fogB4yjP/BHbk4sxDyOCHbNlpCOXR5QoWLzeDK76jTDlowvICawYPVGoikiyS0woGth3okZhREdOISQt99bLWACtua8thk/b/PHxwKA+2MacHXsL3a
fKMGFXmaoogdI3SFTIIveRcuOIc7bqDU6se+IGk74E2rU6TmY4DJMH/U7jpQ6ucV37lUh6u5qRICI4Rv7g/I/sQ1FWCqcP9UCO5rGb6k6GMI5D2ioHIRY1lmSdyuczSp
dPC7WSQQi9M7bkEPm/5NUe3wt9II4iUcSZ39U5N1icRinUdNfitP9jRh2Ps7eCuQFxhF6nLoBjuRYACIgl+aDXTwu1kkEIvTO25BD5v+TVECLKdCJGHP5fs+ax1XOqAY
99MSJRZxm4DhiCBpdeGI5ePlbxnuq7WINR5kEANQ7ALx+ofJhyks9QeSTHmLZG6V5CjSbld7LLOOAjeKzJn/NOrnu/rJUIpudFkjixWvRhmeSLI1n8jZk2FaAGHZka3g
HUl9cZ4CU7KufOxVc7kLRnPZKJHBC/FQFuwMuZPepD0HEspf2EOkUSAJmyprLvRThjs3CtKp57FOOxQ3DyXJ3V228Z44dZe2QbeSyXNCPI5edhlifoyOwtAQVo2srnn5
c2Ze+61A0TRlZx2P03oDPCrviEENj+QYicA7GDdcpnmsI7xhHof9Lp/ARharcu6fegV6MIBcT0QF6s17mOkfJaxVcV5SPIskUNiBAuF1nKt46BlVvE9kdvukKMGZGLZJ
mxZ/Qhhk4ddwI0CRWj9lmDLBRtb5Ox2zlU25m7pe8Xun2yceC0dPWdbHjB/3evaTKVyRfQK3sZD+aATd3GZNSf73+pVA/PF87F4OsbCNj92tSnn5MHw4QPOYVSKLlFrM
yTqBfsWivBuZefLF/ZqGl9ovNhzRhnlVsHxkDt5jcd5yF2BQrTMWjMy1CQKsz5PHF7GPof+J7AdGIgSR18tAH8pJQKOps7zjYiZp0TnOXW7W/9keLqYs6XpdyFOlU42t
0UNptLc6tSqOKk94cnEX3D5+/uStayjc0uWse0YEnwZ5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t6Namz7jcTxeu5U82lcos45
US09kFLzNhnTQgSW4Fo2XCOS1dxmtwgS+GTXHNTfLxJZrGexMORFTq9+vlyE2xbUkzU+DjiSgktTCWS+RI2UdXn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
ef3risZHFCz9C03WU4Hq3jt53sMzKlvUrR1mL38FexYO9WNtsnTwQKxRXPqJZL58gc7oe9fRS1H6Mh4dG9neL3+gnk8rZfGYmULgvToqlaXPmnPpRWswHdZFeRgZ2/Nb
0864bikiUZ0HC2JEx8iX0e3rwZE/sesGvS2rf4KeWoTapjI4znkxO+ldkLQYNJKrlnnX7C0D/sIR9lC7/38Cbn1Hao9JAS8BPjI/7ZrVdneDQsb4Zf4OPXJWY7LMsAgJ
cfPBCJj04ieE/ACPoio3RW8054C5s9kYG+OXOU2cv18o/rBya39HfUv0QP+FXiE+5r3JM5ZSJY5rpjfDP63oPQFk2UCtzmVaCPPNFOFKhqkXmfAMJK6WQE8q28LqWXMD
gNCgwONXm2mJzlJ4BwUFRk4eP8WOK1XiBEBxirS0cMo+O5s11MDBpp77azchU7mQHCCA/Z6qTOf7Zp4fUX7NxiopLM819M1TQMz/mQUcuqC8xVHbZ07BlecEaY3ElJLs
gvIaOn6rkcjiA/VW2sxaqzvZNlNcT2flV8bm1bEbgLR5/euKxkcULP0LTdZTgereef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t5NNt6F0z3DpKOxrf/dvfrf
nnTVuzfcHzEFt96/u4AD0UMtFjYhn0DJRl/y2h0gkVmLrVwWF28+PqNEFnEbW+JWef3risZHFCz9C03WU4Hq3nn964rGRxQs/QtN1lOB6t55/euKxkcULP0LTdZTgere
O3newzMqW9StHWYvfwV7Fg71Y22ydPBArFFc+olkvnyBzuh719FLUfoyHh0b2d4vGq3i81nGygkan2jD335VC3UNtjlhERNDxfuGvFNkvm+oMkt9NFF95pCRlvKzcLTC
fUdqj0kBLwE+Mj/tmtV2dwbujuSoWil6V30k8bhXtV2zXv/M/jXvWwURizm4Ksn9JZMCI7QyxqYXoavezOAj2zPmkZWa+QGRcEEp8OcMlSNNjjhwCCiTZLB1pUaRuaIw
ewcqrDHbNUK3P2UH6rZI9GLkmVql42+zIRnaJOcYrVRyrJdlCIj8oCwRbVXAx9nWHSFUPiBo4BcnJBmXGKLdqr1T6D1ag/U07QgxCX9STdj5wExzkQOg5Ok6Kq6qm9vB
`pragma protect end_protected

endmodule
