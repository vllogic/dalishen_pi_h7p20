// ============================================================
// File Name: rx_dpram_768x32_ahb.v
// IP core  : ethernet_mac_v2 
// Function : RX memory management
// ============================================================

module cme_ip_rx_dpram_768x32_ahb_v3(
        clkw,
        cew,
        aw,
        dw,

        clkr,
        cer,
        ar,
        qr
        );
//protect_encode_begin
`pragma protect begin_protected
`pragma protect version=1
`pragma protect data_block
joqvu!!!dmls<joqvu!!!dfs<joqvu!!!\:;1^!bs<pvuqvu!!\42;1^!rs<!!!!joqvu!!!dmlx<joqvu!!!dfx<joqvu!!!\:;1^!!!bx<joqvu!!!\42;1^!!ex<xjsf!\42;1^!rs`1<xjsf!\42;1^!rs`2<xjsf!\42;1^!rs`3<xjsf!!!!!!!!dfx`1<xjsf!!!!!!!!dfx`2<xjsf!!!!!!!!dfx`3<xjsf!!!!!!!!dfs`1<xjsf!!!!!!!!dfs`2<xjsf!!!!!!!!dfs`3<sfh!!\2;1^!!bs`t<bmxbzt!A!)qptfehf!dmls*!cfhjo!!!bs`t!=>!bs\:;9^<foebttjho!rs!>!)bs`t!>>!3(i1*!@!rs`1!;!!!!!!!!!!!!)bs`t!>>!3(i2*!@!rs`2!;!!!!!!!!!!!!rs`3<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s1`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`1*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`1*-
!/rs)rs`1\42;27^*!!!!*<bttjho!dfx`1!>!dfx!'!)bx\:;9^!>>!3(c1*<bttjho!dfs`1!>!dfs!'!)bs\:;9^!>>!3(c1*<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s1`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`1*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`1*-
!/rs)rs`1\26;1^*!!!!*<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s2`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`2*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`2*-
!/rs)rs`2\42;27^*!!!!*<
!bttjho!dfx`2!>!dfx!'!)bx\:;9^!>>!3(c2*<
bttjho!dfs`2!>!dfs!'!)bs\:;9^!>>!3(c2*<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s2`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`2*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`2*-
!/rs)rs`2\26;1^*!!!!*<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s3`w2)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`3*-
!/ex)ex\42;27^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`3*-
!/rs)rs`3\42;27^*!!!!*<
!bttjho!dfx`3!>!dfx!'!)bx\:;9^!>>!3(c21*<bttjho!dfs`3!>!dfs!'!)bs\:;9^!>>!3(c21*<dnf`jq`fnc6l`fui`n8`w4!fnc`jotu`s3`w1)
!/dmlx)dmlx*-
!/bx)bx\8;1^*-
!/dfx)dfx`3*-
!/ex)ex\26;1^*-

!/dmls)dmls*-
!/bs)bs\8;1^*-
!/dfs)dfs`3*-
!/rs)rs`3\26;1^*!!!!*<
`pragma protect end_protected
//protect_encode_end
endmodule


